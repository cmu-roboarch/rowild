/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_pointsOverlap_double_2 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    axis_address0,
    axis_ce0,
    axis_q0,
    axis_address1,
    axis_ce1,
    axis_q1,
    axis_offset1,
    ap_return
);

    parameter ap_ST_fsm_pp0_stage0 = 14'd1;
    parameter ap_ST_fsm_pp0_stage1 = 14'd2;
    parameter ap_ST_fsm_pp0_stage2 = 14'd4;
    parameter ap_ST_fsm_pp0_stage3 = 14'd8;
    parameter ap_ST_fsm_pp0_stage4 = 14'd16;
    parameter ap_ST_fsm_pp0_stage5 = 14'd32;
    parameter ap_ST_fsm_pp0_stage6 = 14'd64;
    parameter ap_ST_fsm_pp0_stage7 = 14'd128;
    parameter ap_ST_fsm_pp0_stage8 = 14'd256;
    parameter ap_ST_fsm_pp0_stage9 = 14'd512;
    parameter ap_ST_fsm_pp0_stage10 = 14'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 14'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 14'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 14'd8192;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    output [5:0] axis_address0;
    output axis_ce0;
    input [63:0] axis_q0;
    output [5:0] axis_address1;
    output axis_ce1;
    input [63:0] axis_q1;
    input [1:0] axis_offset1;
    output [0:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[6:0] p1_address0;
    reg p1_ce0;
    reg[6:0] p1_address1;
    reg p1_ce1;
    reg p2_0_0_ce0;
    reg p2_0_1_ce0;
    reg p2_0_2_ce0;
    reg p2_1_0_ce0;
    reg p2_1_1_ce0;
    reg p2_1_2_ce0;
    reg p2_2_0_ce0;
    reg p2_2_1_ce0;
    reg p2_2_2_ce0;
    reg p2_3_0_ce0;
    reg p2_3_1_ce0;
    reg p2_3_2_ce0;
    reg p2_4_0_ce0;
    reg p2_4_1_ce0;
    reg p2_4_2_ce0;
    reg p2_5_0_ce0;
    reg p2_5_1_ce0;
    reg p2_5_2_ce0;
    reg p2_6_0_ce0;
    reg p2_6_1_ce0;
    reg p2_6_2_ce0;
    reg p2_7_0_ce0;
    reg p2_7_1_ce0;
    reg p2_7_2_ce0;
    reg p2_8_0_ce0;
    reg p2_8_1_ce0;
    reg p2_8_2_ce0;
    reg[5:0] axis_address0;
    reg axis_ce0;
    reg axis_ce1;

    (* fsm_encoding = "none" *) reg   [13:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_subdone;
    reg   [63:0] reg_819;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    reg   [63:0] reg_824;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    reg   [63:0] reg_830;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    reg   [63:0] reg_835;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    reg   [63:0] reg_842;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    wire    ap_block_pp0_stage13_11001;
    reg   [63:0] reg_849;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] grp_fu_781_p2;
    reg   [63:0] reg_855;
    wire   [63:0] grp_fu_786_p2;
    reg   [63:0] reg_862;
    reg   [63:0] reg_869;
    reg   [63:0] reg_876;
    reg   [63:0] reg_883;
    reg   [63:0] reg_890;
    reg   [63:0] reg_898;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    reg   [63:0] reg_905;
    reg   [63:0] reg_911;
    reg   [63:0] reg_917;
    wire   [63:0] grp_fu_771_p2;
    reg   [63:0] reg_923;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire   [63:0] p2_offset_cast_fu_934_p1;
    reg   [63:0] p2_offset_cast_reg_3746;
    wire   [6:0] mul_ln120_fu_972_p2;
    reg   [6:0] mul_ln120_reg_3751;
    wire   [5:0] add_ln120_2_fu_1005_p2;
    reg   [5:0] add_ln120_2_reg_3786;
    wire   [5:0] sub_ln120_1_fu_1036_p2;
    reg   [5:0] sub_ln120_1_reg_3932;
    reg   [63:0] p1_load_reg_3947;
    reg   [63:0] p2_0_0_load_reg_3952;
    reg   [63:0] p2_0_1_load_reg_3957;
    reg   [63:0] p2_0_2_load_reg_3962;
    reg   [63:0] p2_1_0_load_reg_3967;
    reg   [63:0] p2_1_1_load_reg_3972;
    reg   [63:0] p2_1_2_load_reg_3977;
    reg   [63:0] p2_2_0_load_reg_3982;
    reg   [63:0] p2_2_1_load_reg_3987;
    reg   [63:0] p2_2_2_load_reg_3992;
    reg   [63:0] p2_3_0_load_reg_3997;
    reg   [63:0] p2_3_1_load_reg_4002;
    reg   [63:0] p2_3_2_load_reg_4007;
    reg   [63:0] p2_4_0_load_reg_4012;
    reg   [63:0] p2_4_1_load_reg_4017;
    reg   [63:0] p2_4_2_load_reg_4022;
    reg   [63:0] p2_5_0_load_reg_4027;
    reg   [63:0] p2_5_1_load_reg_4032;
    reg   [63:0] p2_5_2_load_reg_4037;
    reg   [63:0] p2_6_0_load_reg_4042;
    reg   [63:0] p2_6_1_load_reg_4047;
    reg   [63:0] p2_6_2_load_reg_4052;
    reg   [63:0] p2_7_0_load_reg_4057;
    reg   [63:0] p2_7_1_load_reg_4062;
    reg   [63:0] p2_7_2_load_reg_4067;
    reg   [63:0] p2_8_0_load_reg_4072;
    reg   [63:0] p2_8_1_load_reg_4077;
    reg   [63:0] axis_load_reg_4097;
    reg   [63:0] axis_load_1_reg_4105;
    reg   [63:0] p1_load_6_reg_4113;
    reg   [63:0] axis_load_2_reg_4128;
    reg   [63:0] p1_load_12_reg_4136;
    reg   [63:0] p1_load_4_reg_4151;
    reg   [63:0] p1_load_7_reg_4166;
    reg   [63:0] p1_load_10_reg_4181;
    reg   [63:0] p1_load_13_reg_4196;
    reg   [63:0] p1_load_2_reg_4211;
    reg   [63:0] p1_load_5_reg_4216;
    wire   [63:0] grp_fu_791_p2;
    reg   [63:0] mul_reg_4231;
    wire   [63:0] grp_fu_795_p2;
    reg   [63:0] mul6_reg_4236;
    wire   [63:0] grp_fu_799_p2;
    reg   [63:0] mul1_reg_4241;
    wire   [63:0] grp_fu_803_p2;
    reg   [63:0] mul2_reg_4246;
    reg   [63:0] p1_load_16_reg_4251;
    reg   [63:0] mul20_1_reg_4266;
    reg   [63:0] mul25_1_reg_4271;
    reg   [63:0] mul20_2_reg_4276;
    reg   [63:0] mul25_2_reg_4281;
    reg   [63:0] p1_load_19_reg_4286;
    reg   [63:0] mul_1_reg_4301;
    reg   [63:0] mul6_1_reg_4306;
    reg   [63:0] mul20_3_reg_4311;
    reg   [63:0] mul25_3_reg_4316;
    reg   [63:0] p1_load_22_reg_4321;
    reg   [63:0] mul20_s_reg_4336;
    reg   [63:0] mul25_s_reg_4341;
    reg   [63:0] mul20_4_reg_4346;
    reg   [63:0] mul25_4_reg_4351;
    reg   [63:0] p1_load_25_reg_4356;
    reg   [63:0] mul20_1_1_reg_4371;
    reg   [63:0] mul25_1_1_reg_4376;
    reg   [63:0] mul20_5_reg_4381;
    reg   [63:0] mul25_5_reg_4386;
    reg   [63:0] p1_load_20_reg_4391;
    reg   [63:0] mul20_2_1_reg_4396;
    reg   [63:0] mul25_2_1_reg_4401;
    reg   [63:0] mul20_6_reg_4406;
    reg   [63:0] mul25_6_reg_4411;
    reg   [63:0] p1_load_26_reg_4416;
    reg   [63:0] mul_2_reg_4426;
    reg   [63:0] mul6_2_reg_4431;
    reg   [63:0] mul20_3_1_reg_4436;
    reg   [63:0] mul25_3_1_reg_4441;
    reg   [63:0] p2_8_2_load_reg_4446;
    reg   [63:0] max1_11_reg_4451;
    wire   [63:0] grp_fu_776_p2;
    reg   [63:0] max2_11_reg_4456;
    reg   [63:0] mul20_8_reg_4461;
    reg   [63:0] mul25_8_reg_4466;
    reg   [63:0] mul20_7_reg_4471;
    reg   [63:0] mul25_7_reg_4476;
    reg   [63:0] n1_3_reg_4481;
    reg   [63:0] n2_3_reg_4486;
    reg   [63:0] mul20_1_2_reg_4491;
    reg   [63:0] mul25_1_2_reg_4496;
    reg   [63:0] n2_6_reg_4501;
    reg   [63:0] mul20_4_1_reg_4506;
    reg   [63:0] mul25_4_1_reg_4511;
    reg   [63:0] mul20_2_2_reg_4516;
    reg   [63:0] mul25_2_2_reg_4521;
    reg   [63:0] n1_9_reg_4526;
    reg   [63:0] n2_9_reg_4531;
    reg   [63:0] mul20_5_1_reg_4536;
    reg   [63:0] mul25_5_1_reg_4541;
    reg   [63:0] mul20_3_2_reg_4546;
    reg   [63:0] mul25_3_2_reg_4551;
    reg   [63:0] n1_12_reg_4556;
    reg   [63:0] n2_12_reg_4561;
    reg   [63:0] mul20_6_1_reg_4566;
    reg   [63:0] mul25_6_1_reg_4571;
    reg   [63:0] mul20_4_2_reg_4576;
    reg   [63:0] mul25_4_2_reg_4581;
    reg   [63:0] n1_15_reg_4586;
    reg   [63:0] n2_15_reg_4591;
    reg   [63:0] mul20_7_1_reg_4596;
    reg   [63:0] mul25_7_1_reg_4601;
    reg   [63:0] mul20_5_2_reg_4606;
    reg   [63:0] mul25_5_2_reg_4611;
    reg   [63:0] n1_18_reg_4616;
    reg   [63:0] n2_18_reg_4621;
    reg   [63:0] mul20_6_2_reg_4626;
    reg   [63:0] mul20_6_2_reg_4626_pp0_iter2_reg;
    reg   [63:0] mul25_6_2_reg_4631;
    reg   [63:0] mul25_6_2_reg_4631_pp0_iter2_reg;
    reg   [63:0] mul20_7_2_reg_4636;
    reg   [63:0] mul20_7_2_reg_4636_pp0_iter2_reg;
    reg   [63:0] mul25_7_2_reg_4641;
    reg   [63:0] mul25_7_2_reg_4641_pp0_iter2_reg;
    reg   [63:0] max1_1_reg_4646;
    reg   [63:0] max2_1_reg_4651;
    reg   [63:0] n1_4_reg_4656;
    reg   [63:0] n2_4_reg_4661;
    reg   [63:0] n1_7_reg_4666;
    reg   [63:0] n2_7_reg_4671;
    reg   [63:0] n1_10_reg_4676;
    reg   [63:0] n2_10_reg_4681;
    reg   [63:0] n1_21_reg_4686;
    reg   [63:0] n2_21_reg_4691;
    reg   [63:0] n1_13_reg_4696;
    reg   [63:0] n2_13_reg_4701;
    reg   [63:0] n1_16_reg_4706;
    reg   [63:0] n2_16_reg_4711;
    reg   [63:0] n1_19_reg_4716;
    reg   [63:0] n2_19_reg_4721;
    wire   [63:0] max1_fu_1391_p3;
    reg   [63:0] max1_reg_4726;
    wire   [63:0] min1_2_fu_1405_p3;
    reg   [63:0] min1_2_reg_4733;
    wire   [0:0] and_ln135_fu_1485_p2;
    reg   [0:0] and_ln135_reg_4740;
    wire   [0:0] grp_fu_815_p2;
    reg   [0:0] tmp_9_reg_4746;
    wire   [63:0] max2_fu_1495_p3;
    reg   [63:0] max2_reg_4751;
    wire   [63:0] min2_2_fu_1509_p3;
    reg   [63:0] min2_2_reg_4758;
    reg   [63:0] n2_11_reg_4765;
    reg   [63:0] n1_22_reg_4774;
    wire   [63:0] max1_4_fu_1600_p3;
    reg   [63:0] max1_4_reg_4779;
    wire   [63:0] min1_3_fu_1654_p3;
    reg   [63:0] min1_3_reg_4786;
    wire   [0:0] or_ln135_2_fu_1708_p2;
    reg   [0:0] or_ln135_2_reg_4793;
    wire   [63:0] max2_4_fu_1744_p3;
    reg   [63:0] max2_4_reg_4798;
    wire   [63:0] min2_3_fu_1797_p3;
    reg   [63:0] min2_3_reg_4805;
    wire   [63:0] max1_5_fu_1887_p3;
    reg   [63:0] max1_5_reg_4812;
    wire   [63:0] min1_4_fu_1941_p3;
    reg   [63:0] min1_4_reg_4819;
    wire   [0:0] or_ln135_4_fu_1995_p2;
    reg   [0:0] or_ln135_4_reg_4826;
    wire   [63:0] max2_5_fu_2031_p3;
    reg   [63:0] max2_5_reg_4831;
    wire   [63:0] min2_4_fu_2084_p3;
    reg   [63:0] min2_4_reg_4838;
    wire   [63:0] max1_6_fu_2174_p3;
    reg   [63:0] max1_6_reg_4845;
    wire   [63:0] min1_5_fu_2228_p3;
    reg   [63:0] min1_5_reg_4852;
    wire   [0:0] or_ln135_6_fu_2281_p2;
    reg   [0:0] or_ln135_6_reg_4859;
    wire   [63:0] max2_6_fu_2317_p3;
    reg   [63:0] max2_6_reg_4864;
    wire   [63:0] min2_5_fu_2369_p3;
    reg   [63:0] min2_5_reg_4871;
    wire   [63:0] max1_7_fu_2458_p3;
    reg   [63:0] max1_7_reg_4878;
    wire   [63:0] min1_6_fu_2512_p3;
    reg   [63:0] min1_6_reg_4885;
    wire   [0:0] or_ln135_8_fu_2566_p2;
    reg   [0:0] or_ln135_8_reg_4892;
    wire   [63:0] max2_7_fu_2602_p3;
    reg   [63:0] max2_7_reg_4897;
    reg   [63:0] n2_23_reg_4904;
    wire   [63:0] min2_6_fu_2655_p3;
    reg   [63:0] min2_6_reg_4913;
    wire   [63:0] max1_8_fu_2745_p3;
    reg   [63:0] max1_8_reg_4920;
    wire   [63:0] min1_7_fu_2799_p3;
    reg   [63:0] min1_7_reg_4927;
    wire   [0:0] or_ln135_10_fu_2853_p2;
    reg   [0:0] or_ln135_10_reg_4934;
    wire   [63:0] max2_8_fu_2889_p3;
    reg   [63:0] max2_8_reg_4939;
    wire   [63:0] min2_7_fu_2942_p3;
    reg   [63:0] min2_7_reg_4946;
    wire   [63:0] max1_9_fu_3032_p3;
    reg   [63:0] max1_9_reg_4953;
    wire   [63:0] min1_8_fu_3086_p3;
    reg   [63:0] min1_8_reg_4960;
    wire   [0:0] or_ln135_12_fu_3140_p2;
    reg   [0:0] or_ln135_12_reg_4967;
    wire   [63:0] max2_9_fu_3176_p3;
    reg   [63:0] max2_9_reg_4972;
    wire   [63:0] min2_8_fu_3229_p3;
    reg   [63:0] min2_8_reg_4979;
    wire   [63:0] max1_10_fu_3319_p3;
    reg   [63:0] max1_10_reg_4986;
    wire   [63:0] min1_9_fu_3373_p3;
    reg   [63:0] min1_9_reg_4993;
    wire   [63:0] max2_10_fu_3462_p3;
    reg   [63:0] max2_10_reg_5001;
    wire   [63:0] min2_9_fu_3515_p3;
    reg   [63:0] min2_9_reg_5009;
    wire   [0:0] grp_fu_811_p2;
    reg   [0:0] tmp_82_reg_5016;
    reg   [0:0] tmp_84_reg_5021;
    reg   [0:0] tmp_85_reg_5026;
    reg   [0:0] tmp_86_reg_5031;
    wire   [0:0] and_ln139_1_fu_3591_p2;
    reg   [0:0] and_ln139_1_reg_5036;
    wire   [0:0] and_ln139_4_fu_3638_p2;
    reg   [0:0] and_ln139_4_reg_5041;
    wire   [0:0] and_ln140_3_fu_3689_p2;
    reg   [0:0] and_ln140_3_reg_5047;
    wire   [0:0] and_ln140_fu_3711_p2;
    reg   [0:0] and_ln140_reg_5052;
    reg   [0:0] tmp_80_reg_5057;
    wire   [0:0] or_ln140_2_fu_3727_p2;
    reg   [0:0] or_ln140_2_reg_5062;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage3_subdone;
    wire   [63:0] zext_ln120_2_fu_978_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln129_fu_1016_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln129_3_fu_1026_p1;
    wire   [63:0] zext_ln120_6_fu_1041_p1;
    wire   [63:0] zext_ln120_7_fu_1052_p1;
    wire   [63:0] zext_ln129_6_fu_1062_p1;
    wire    ap_block_pp0_stage2;
    wire   [63:0] zext_ln129_9_fu_1072_p1;
    wire   [63:0] zext_ln120_8_fu_1082_p1;
    wire   [63:0] zext_ln120_3_fu_1092_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln129_1_fu_1102_p1;
    wire   [63:0] zext_ln129_4_fu_1112_p1;
    wire    ap_block_pp0_stage4;
    wire   [63:0] zext_ln129_12_fu_1122_p1;
    wire   [63:0] zext_ln129_7_fu_1132_p1;
    wire    ap_block_pp0_stage5;
    wire   [63:0] zext_ln129_15_fu_1142_p1;
    wire   [63:0] zext_ln129_10_fu_1152_p1;
    wire    ap_block_pp0_stage6;
    wire   [63:0] zext_ln129_18_fu_1162_p1;
    wire   [63:0] zext_ln120_4_fu_1172_p1;
    wire    ap_block_pp0_stage7;
    wire   [63:0] zext_ln129_2_fu_1182_p1;
    wire   [63:0] zext_ln129_13_fu_1192_p1;
    wire    ap_block_pp0_stage8;
    wire   [63:0] zext_ln129_21_fu_1202_p1;
    wire   [63:0] zext_ln129_5_fu_1212_p1;
    wire    ap_block_pp0_stage9;
    wire   [63:0] zext_ln129_16_fu_1222_p1;
    wire   [63:0] zext_ln129_8_fu_1232_p1;
    wire    ap_block_pp0_stage10;
    wire   [63:0] zext_ln129_19_fu_1242_p1;
    wire   [63:0] zext_ln129_11_fu_1252_p1;
    wire    ap_block_pp0_stage11;
    wire   [63:0] zext_ln129_22_fu_1262_p1;
    wire   [63:0] zext_ln129_14_fu_1272_p1;
    wire    ap_block_pp0_stage12;
    wire   [63:0] zext_ln129_17_fu_1282_p1;
    wire   [63:0] zext_ln129_20_fu_1292_p1;
    wire    ap_block_pp0_stage13;
    wire   [63:0] zext_ln129_23_fu_1302_p1;
    reg   [63:0] grp_fu_771_p0;
    reg   [63:0] grp_fu_771_p1;
    reg   [63:0] grp_fu_776_p0;
    reg   [63:0] grp_fu_776_p1;
    reg   [63:0] grp_fu_781_p0;
    reg   [63:0] grp_fu_781_p1;
    reg   [63:0] grp_fu_786_p0;
    reg   [63:0] grp_fu_786_p1;
    reg   [63:0] grp_fu_791_p0;
    reg   [63:0] grp_fu_791_p1;
    reg   [63:0] grp_fu_795_p0;
    reg   [63:0] grp_fu_795_p1;
    reg   [63:0] grp_fu_799_p0;
    reg   [63:0] grp_fu_799_p1;
    reg   [63:0] grp_fu_803_p0;
    reg   [63:0] grp_fu_803_p1;
    reg   [63:0] grp_fu_807_p0;
    reg   [63:0] grp_fu_807_p1;
    reg   [63:0] grp_fu_811_p0;
    reg   [63:0] grp_fu_811_p1;
    reg   [63:0] grp_fu_815_p0;
    reg   [63:0] grp_fu_815_p1;
    wire   [1:0] mul_ln120_fu_972_p0;
    wire   [5:0] mul_ln120_fu_972_p1;
    wire   [3:0] tmp_fu_983_p3;
    wire   [4:0] zext_ln120_5_fu_991_p1;
    wire   [4:0] zext_ln120_fu_964_p1;
    wire   [4:0] sub_ln120_fu_995_p2;
    wire  signed [5:0] sext_ln120_fu_1001_p1;
    wire   [5:0] axis_offset1_cast4_fu_930_p1;
    wire   [6:0] add_ln129_fu_1011_p2;
    wire   [6:0] add_ln129_3_fu_1021_p2;
    wire   [5:0] shl_ln120_fu_1031_p2;
    wire   [5:0] add_ln120_3_fu_1046_p2;
    wire   [6:0] add_ln129_6_fu_1057_p2;
    wire   [6:0] add_ln129_9_fu_1067_p2;
    wire   [5:0] add_ln120_4_fu_1077_p2;
    wire   [6:0] add_ln120_fu_1087_p2;
    wire   [6:0] add_ln129_1_fu_1097_p2;
    wire   [6:0] add_ln129_4_fu_1107_p2;
    wire   [6:0] add_ln129_12_fu_1117_p2;
    wire   [6:0] add_ln129_7_fu_1127_p2;
    wire   [6:0] add_ln129_15_fu_1137_p2;
    wire   [6:0] add_ln129_10_fu_1147_p2;
    wire   [6:0] add_ln129_18_fu_1157_p2;
    wire   [6:0] add_ln120_1_fu_1167_p2;
    wire   [6:0] add_ln129_2_fu_1177_p2;
    wire   [6:0] add_ln129_13_fu_1187_p2;
    wire   [6:0] add_ln129_21_fu_1197_p2;
    wire   [6:0] add_ln129_5_fu_1207_p2;
    wire   [6:0] add_ln129_16_fu_1217_p2;
    wire   [6:0] add_ln129_8_fu_1227_p2;
    wire   [6:0] add_ln129_19_fu_1237_p2;
    wire   [6:0] add_ln129_11_fu_1247_p2;
    wire   [6:0] add_ln129_22_fu_1257_p2;
    wire   [6:0] add_ln129_14_fu_1267_p2;
    wire   [6:0] add_ln129_17_fu_1277_p2;
    wire   [6:0] add_ln129_20_fu_1287_p2;
    wire   [6:0] add_ln129_23_fu_1297_p2;
    wire   [63:0] bitcast_ln133_fu_1307_p1;
    wire   [63:0] bitcast_ln133_1_fu_1325_p1;
    wire   [10:0] tmp_1_fu_1311_p4;
    wire   [51:0] trunc_ln133_fu_1321_p1;
    wire   [0:0] icmp_ln133_1_fu_1349_p2;
    wire   [0:0] icmp_ln133_fu_1343_p2;
    wire   [10:0] tmp_2_fu_1329_p4;
    wire   [51:0] trunc_ln133_1_fu_1339_p1;
    wire   [0:0] icmp_ln133_3_fu_1367_p2;
    wire   [0:0] icmp_ln133_2_fu_1361_p2;
    wire   [0:0] or_ln133_fu_1355_p2;
    wire   [0:0] or_ln133_1_fu_1373_p2;
    wire   [0:0] and_ln133_fu_1379_p2;
    wire   [0:0] grp_fu_807_p2;
    wire   [0:0] and_ln133_1_fu_1385_p2;
    wire   [0:0] and_ln134_fu_1399_p2;
    wire   [63:0] bitcast_ln135_fu_1413_p1;
    wire   [63:0] bitcast_ln135_1_fu_1431_p1;
    wire   [10:0] tmp_7_fu_1417_p4;
    wire   [51:0] trunc_ln135_fu_1427_p1;
    wire   [0:0] icmp_ln135_1_fu_1455_p2;
    wire   [0:0] icmp_ln135_fu_1449_p2;
    wire   [10:0] tmp_8_fu_1435_p4;
    wire   [51:0] trunc_ln135_1_fu_1445_p1;
    wire   [0:0] icmp_ln135_3_fu_1473_p2;
    wire   [0:0] icmp_ln135_2_fu_1467_p2;
    wire   [0:0] or_ln135_fu_1461_p2;
    wire   [0:0] or_ln135_1_fu_1479_p2;
    wire   [0:0] and_ln135_1_fu_1491_p2;
    wire   [0:0] and_ln136_fu_1504_p2;
    wire   [63:0] bitcast_ln133_2_fu_1517_p1;
    wire   [63:0] bitcast_ln133_3_fu_1535_p1;
    wire   [10:0] tmp_4_fu_1521_p4;
    wire   [51:0] trunc_ln133_2_fu_1531_p1;
    wire   [0:0] icmp_ln133_5_fu_1558_p2;
    wire   [0:0] icmp_ln133_4_fu_1552_p2;
    wire   [10:0] tmp_5_fu_1538_p4;
    wire   [51:0] trunc_ln133_3_fu_1548_p1;
    wire   [0:0] icmp_ln133_7_fu_1576_p2;
    wire   [0:0] icmp_ln133_6_fu_1570_p2;
    wire   [0:0] or_ln133_2_fu_1564_p2;
    wire   [0:0] or_ln133_3_fu_1582_p2;
    wire   [0:0] and_ln133_2_fu_1588_p2;
    wire   [0:0] and_ln133_3_fu_1594_p2;
    wire   [63:0] bitcast_ln134_fu_1607_p1;
    wire   [10:0] tmp_11_fu_1610_p4;
    wire   [51:0] trunc_ln134_fu_1620_p1;
    wire   [0:0] icmp_ln134_1_fu_1630_p2;
    wire   [0:0] icmp_ln134_fu_1624_p2;
    wire   [0:0] or_ln134_fu_1636_p2;
    wire   [0:0] and_ln134_1_fu_1642_p2;
    wire   [0:0] and_ln134_2_fu_1648_p2;
    wire   [63:0] bitcast_ln135_2_fu_1661_p1;
    wire   [63:0] bitcast_ln135_3_fu_1679_p1;
    wire   [10:0] tmp_13_fu_1665_p4;
    wire   [51:0] trunc_ln135_2_fu_1675_p1;
    wire   [0:0] icmp_ln135_5_fu_1702_p2;
    wire   [0:0] icmp_ln135_4_fu_1696_p2;
    wire   [10:0] tmp_14_fu_1682_p4;
    wire   [51:0] trunc_ln135_3_fu_1692_p1;
    wire   [0:0] icmp_ln135_7_fu_1720_p2;
    wire   [0:0] icmp_ln135_6_fu_1714_p2;
    wire   [0:0] or_ln135_3_fu_1726_p2;
    wire   [0:0] and_ln135_2_fu_1732_p2;
    wire   [0:0] and_ln135_3_fu_1738_p2;
    wire   [63:0] bitcast_ln136_fu_1751_p1;
    wire   [10:0] tmp_16_fu_1754_p4;
    wire   [51:0] trunc_ln136_fu_1764_p1;
    wire   [0:0] icmp_ln136_1_fu_1774_p2;
    wire   [0:0] icmp_ln136_fu_1768_p2;
    wire   [0:0] or_ln136_fu_1780_p2;
    wire   [0:0] and_ln136_1_fu_1786_p2;
    wire   [0:0] and_ln136_2_fu_1791_p2;
    wire   [63:0] bitcast_ln133_4_fu_1804_p1;
    wire   [63:0] bitcast_ln133_5_fu_1822_p1;
    wire   [10:0] tmp_18_fu_1808_p4;
    wire   [51:0] trunc_ln133_4_fu_1818_p1;
    wire   [0:0] icmp_ln133_9_fu_1845_p2;
    wire   [0:0] icmp_ln133_8_fu_1839_p2;
    wire   [10:0] tmp_19_fu_1825_p4;
    wire   [51:0] trunc_ln133_5_fu_1835_p1;
    wire   [0:0] icmp_ln133_11_fu_1863_p2;
    wire   [0:0] icmp_ln133_10_fu_1857_p2;
    wire   [0:0] or_ln133_4_fu_1851_p2;
    wire   [0:0] or_ln133_5_fu_1869_p2;
    wire   [0:0] and_ln133_4_fu_1875_p2;
    wire   [0:0] and_ln133_5_fu_1881_p2;
    wire   [63:0] bitcast_ln134_1_fu_1894_p1;
    wire   [10:0] tmp_21_fu_1897_p4;
    wire   [51:0] trunc_ln134_1_fu_1907_p1;
    wire   [0:0] icmp_ln134_3_fu_1917_p2;
    wire   [0:0] icmp_ln134_2_fu_1911_p2;
    wire   [0:0] or_ln134_1_fu_1923_p2;
    wire   [0:0] and_ln134_3_fu_1929_p2;
    wire   [0:0] and_ln134_4_fu_1935_p2;
    wire   [63:0] bitcast_ln135_4_fu_1948_p1;
    wire   [63:0] bitcast_ln135_5_fu_1966_p1;
    wire   [10:0] tmp_23_fu_1952_p4;
    wire   [51:0] trunc_ln135_4_fu_1962_p1;
    wire   [0:0] icmp_ln135_9_fu_1989_p2;
    wire   [0:0] icmp_ln135_8_fu_1983_p2;
    wire   [10:0] tmp_24_fu_1969_p4;
    wire   [51:0] trunc_ln135_5_fu_1979_p1;
    wire   [0:0] icmp_ln135_11_fu_2007_p2;
    wire   [0:0] icmp_ln135_10_fu_2001_p2;
    wire   [0:0] or_ln135_5_fu_2013_p2;
    wire   [0:0] and_ln135_4_fu_2019_p2;
    wire   [0:0] and_ln135_5_fu_2025_p2;
    wire   [63:0] bitcast_ln136_1_fu_2038_p1;
    wire   [10:0] tmp_26_fu_2041_p4;
    wire   [51:0] trunc_ln136_1_fu_2051_p1;
    wire   [0:0] icmp_ln136_3_fu_2061_p2;
    wire   [0:0] icmp_ln136_2_fu_2055_p2;
    wire   [0:0] or_ln136_1_fu_2067_p2;
    wire   [0:0] and_ln136_3_fu_2073_p2;
    wire   [0:0] and_ln136_4_fu_2078_p2;
    wire   [63:0] bitcast_ln133_6_fu_2091_p1;
    wire   [63:0] bitcast_ln133_7_fu_2109_p1;
    wire   [10:0] tmp_28_fu_2095_p4;
    wire   [51:0] trunc_ln133_6_fu_2105_p1;
    wire   [0:0] icmp_ln133_13_fu_2132_p2;
    wire   [0:0] icmp_ln133_12_fu_2126_p2;
    wire   [10:0] tmp_29_fu_2112_p4;
    wire   [51:0] trunc_ln133_7_fu_2122_p1;
    wire   [0:0] icmp_ln133_15_fu_2150_p2;
    wire   [0:0] icmp_ln133_14_fu_2144_p2;
    wire   [0:0] or_ln133_6_fu_2138_p2;
    wire   [0:0] or_ln133_7_fu_2156_p2;
    wire   [0:0] and_ln133_6_fu_2162_p2;
    wire   [0:0] and_ln133_7_fu_2168_p2;
    wire   [63:0] bitcast_ln134_2_fu_2181_p1;
    wire   [10:0] tmp_31_fu_2184_p4;
    wire   [51:0] trunc_ln134_2_fu_2194_p1;
    wire   [0:0] icmp_ln134_5_fu_2204_p2;
    wire   [0:0] icmp_ln134_4_fu_2198_p2;
    wire   [0:0] or_ln134_2_fu_2210_p2;
    wire   [0:0] and_ln134_5_fu_2216_p2;
    wire   [0:0] and_ln134_6_fu_2222_p2;
    wire   [63:0] bitcast_ln135_6_fu_2235_p1;
    wire   [63:0] bitcast_ln135_7_fu_2252_p1;
    wire   [10:0] tmp_33_fu_2238_p4;
    wire   [51:0] trunc_ln135_6_fu_2248_p1;
    wire   [0:0] icmp_ln135_13_fu_2275_p2;
    wire   [0:0] icmp_ln135_12_fu_2269_p2;
    wire   [10:0] tmp_34_fu_2255_p4;
    wire   [51:0] trunc_ln135_7_fu_2265_p1;
    wire   [0:0] icmp_ln135_15_fu_2293_p2;
    wire   [0:0] icmp_ln135_14_fu_2287_p2;
    wire   [0:0] or_ln135_7_fu_2299_p2;
    wire   [0:0] and_ln135_6_fu_2305_p2;
    wire   [0:0] and_ln135_7_fu_2311_p2;
    wire   [63:0] bitcast_ln136_2_fu_2323_p1;
    wire   [10:0] tmp_36_fu_2326_p4;
    wire   [51:0] trunc_ln136_2_fu_2336_p1;
    wire   [0:0] icmp_ln136_5_fu_2346_p2;
    wire   [0:0] icmp_ln136_4_fu_2340_p2;
    wire   [0:0] or_ln136_2_fu_2352_p2;
    wire   [0:0] and_ln136_5_fu_2358_p2;
    wire   [0:0] and_ln136_6_fu_2363_p2;
    wire   [63:0] bitcast_ln133_8_fu_2375_p1;
    wire   [63:0] bitcast_ln133_9_fu_2393_p1;
    wire   [10:0] tmp_38_fu_2379_p4;
    wire   [51:0] trunc_ln133_8_fu_2389_p1;
    wire   [0:0] icmp_ln133_17_fu_2416_p2;
    wire   [0:0] icmp_ln133_16_fu_2410_p2;
    wire   [10:0] tmp_39_fu_2396_p4;
    wire   [51:0] trunc_ln133_9_fu_2406_p1;
    wire   [0:0] icmp_ln133_19_fu_2434_p2;
    wire   [0:0] icmp_ln133_18_fu_2428_p2;
    wire   [0:0] or_ln133_8_fu_2422_p2;
    wire   [0:0] or_ln133_9_fu_2440_p2;
    wire   [0:0] and_ln133_8_fu_2446_p2;
    wire   [0:0] and_ln133_9_fu_2452_p2;
    wire   [63:0] bitcast_ln134_3_fu_2465_p1;
    wire   [10:0] tmp_41_fu_2468_p4;
    wire   [51:0] trunc_ln134_3_fu_2478_p1;
    wire   [0:0] icmp_ln134_7_fu_2488_p2;
    wire   [0:0] icmp_ln134_6_fu_2482_p2;
    wire   [0:0] or_ln134_3_fu_2494_p2;
    wire   [0:0] and_ln134_7_fu_2500_p2;
    wire   [0:0] and_ln134_8_fu_2506_p2;
    wire   [63:0] bitcast_ln135_8_fu_2519_p1;
    wire   [63:0] bitcast_ln135_9_fu_2537_p1;
    wire   [10:0] tmp_43_fu_2523_p4;
    wire   [51:0] trunc_ln135_8_fu_2533_p1;
    wire   [0:0] icmp_ln135_17_fu_2560_p2;
    wire   [0:0] icmp_ln135_16_fu_2554_p2;
    wire   [10:0] tmp_44_fu_2540_p4;
    wire   [51:0] trunc_ln135_9_fu_2550_p1;
    wire   [0:0] icmp_ln135_19_fu_2578_p2;
    wire   [0:0] icmp_ln135_18_fu_2572_p2;
    wire   [0:0] or_ln135_9_fu_2584_p2;
    wire   [0:0] and_ln135_8_fu_2590_p2;
    wire   [0:0] and_ln135_9_fu_2596_p2;
    wire   [63:0] bitcast_ln136_3_fu_2609_p1;
    wire   [10:0] tmp_46_fu_2612_p4;
    wire   [51:0] trunc_ln136_3_fu_2622_p1;
    wire   [0:0] icmp_ln136_7_fu_2632_p2;
    wire   [0:0] icmp_ln136_6_fu_2626_p2;
    wire   [0:0] or_ln136_3_fu_2638_p2;
    wire   [0:0] and_ln136_7_fu_2644_p2;
    wire   [0:0] and_ln136_8_fu_2649_p2;
    wire   [63:0] bitcast_ln133_10_fu_2662_p1;
    wire   [63:0] bitcast_ln133_11_fu_2680_p1;
    wire   [10:0] tmp_48_fu_2666_p4;
    wire   [51:0] trunc_ln133_10_fu_2676_p1;
    wire   [0:0] icmp_ln133_21_fu_2703_p2;
    wire   [0:0] icmp_ln133_20_fu_2697_p2;
    wire   [10:0] tmp_49_fu_2683_p4;
    wire   [51:0] trunc_ln133_11_fu_2693_p1;
    wire   [0:0] icmp_ln133_23_fu_2721_p2;
    wire   [0:0] icmp_ln133_22_fu_2715_p2;
    wire   [0:0] or_ln133_10_fu_2709_p2;
    wire   [0:0] or_ln133_11_fu_2727_p2;
    wire   [0:0] and_ln133_10_fu_2733_p2;
    wire   [0:0] and_ln133_11_fu_2739_p2;
    wire   [63:0] bitcast_ln134_4_fu_2752_p1;
    wire   [10:0] tmp_51_fu_2755_p4;
    wire   [51:0] trunc_ln134_4_fu_2765_p1;
    wire   [0:0] icmp_ln134_9_fu_2775_p2;
    wire   [0:0] icmp_ln134_8_fu_2769_p2;
    wire   [0:0] or_ln134_4_fu_2781_p2;
    wire   [0:0] and_ln134_9_fu_2787_p2;
    wire   [0:0] and_ln134_10_fu_2793_p2;
    wire   [63:0] bitcast_ln135_10_fu_2806_p1;
    wire   [63:0] bitcast_ln135_11_fu_2824_p1;
    wire   [10:0] tmp_53_fu_2810_p4;
    wire   [51:0] trunc_ln135_10_fu_2820_p1;
    wire   [0:0] icmp_ln135_21_fu_2847_p2;
    wire   [0:0] icmp_ln135_20_fu_2841_p2;
    wire   [10:0] tmp_54_fu_2827_p4;
    wire   [51:0] trunc_ln135_11_fu_2837_p1;
    wire   [0:0] icmp_ln135_23_fu_2865_p2;
    wire   [0:0] icmp_ln135_22_fu_2859_p2;
    wire   [0:0] or_ln135_11_fu_2871_p2;
    wire   [0:0] and_ln135_10_fu_2877_p2;
    wire   [0:0] and_ln135_11_fu_2883_p2;
    wire   [63:0] bitcast_ln136_4_fu_2896_p1;
    wire   [10:0] tmp_56_fu_2899_p4;
    wire   [51:0] trunc_ln136_4_fu_2909_p1;
    wire   [0:0] icmp_ln136_9_fu_2919_p2;
    wire   [0:0] icmp_ln136_8_fu_2913_p2;
    wire   [0:0] or_ln136_4_fu_2925_p2;
    wire   [0:0] and_ln136_9_fu_2931_p2;
    wire   [0:0] and_ln136_10_fu_2936_p2;
    wire   [63:0] bitcast_ln133_12_fu_2949_p1;
    wire   [63:0] bitcast_ln133_13_fu_2967_p1;
    wire   [10:0] tmp_58_fu_2953_p4;
    wire   [51:0] trunc_ln133_12_fu_2963_p1;
    wire   [0:0] icmp_ln133_25_fu_2990_p2;
    wire   [0:0] icmp_ln133_24_fu_2984_p2;
    wire   [10:0] tmp_59_fu_2970_p4;
    wire   [51:0] trunc_ln133_13_fu_2980_p1;
    wire   [0:0] icmp_ln133_27_fu_3008_p2;
    wire   [0:0] icmp_ln133_26_fu_3002_p2;
    wire   [0:0] or_ln133_12_fu_2996_p2;
    wire   [0:0] or_ln133_13_fu_3014_p2;
    wire   [0:0] and_ln133_12_fu_3020_p2;
    wire   [0:0] and_ln133_13_fu_3026_p2;
    wire   [63:0] bitcast_ln134_5_fu_3039_p1;
    wire   [10:0] tmp_61_fu_3042_p4;
    wire   [51:0] trunc_ln134_5_fu_3052_p1;
    wire   [0:0] icmp_ln134_11_fu_3062_p2;
    wire   [0:0] icmp_ln134_10_fu_3056_p2;
    wire   [0:0] or_ln134_5_fu_3068_p2;
    wire   [0:0] and_ln134_11_fu_3074_p2;
    wire   [0:0] and_ln134_12_fu_3080_p2;
    wire   [63:0] bitcast_ln135_12_fu_3093_p1;
    wire   [63:0] bitcast_ln135_13_fu_3111_p1;
    wire   [10:0] tmp_63_fu_3097_p4;
    wire   [51:0] trunc_ln135_12_fu_3107_p1;
    wire   [0:0] icmp_ln135_25_fu_3134_p2;
    wire   [0:0] icmp_ln135_24_fu_3128_p2;
    wire   [10:0] tmp_64_fu_3114_p4;
    wire   [51:0] trunc_ln135_13_fu_3124_p1;
    wire   [0:0] icmp_ln135_27_fu_3152_p2;
    wire   [0:0] icmp_ln135_26_fu_3146_p2;
    wire   [0:0] or_ln135_13_fu_3158_p2;
    wire   [0:0] and_ln135_12_fu_3164_p2;
    wire   [0:0] and_ln135_13_fu_3170_p2;
    wire   [63:0] bitcast_ln136_5_fu_3183_p1;
    wire   [10:0] tmp_66_fu_3186_p4;
    wire   [51:0] trunc_ln136_5_fu_3196_p1;
    wire   [0:0] icmp_ln136_11_fu_3206_p2;
    wire   [0:0] icmp_ln136_10_fu_3200_p2;
    wire   [0:0] or_ln136_5_fu_3212_p2;
    wire   [0:0] and_ln136_11_fu_3218_p2;
    wire   [0:0] and_ln136_12_fu_3223_p2;
    wire   [63:0] bitcast_ln133_14_fu_3236_p1;
    wire   [63:0] bitcast_ln133_15_fu_3254_p1;
    wire   [10:0] tmp_68_fu_3240_p4;
    wire   [51:0] trunc_ln133_14_fu_3250_p1;
    wire   [0:0] icmp_ln133_29_fu_3277_p2;
    wire   [0:0] icmp_ln133_28_fu_3271_p2;
    wire   [10:0] tmp_69_fu_3257_p4;
    wire   [51:0] trunc_ln133_15_fu_3267_p1;
    wire   [0:0] icmp_ln133_31_fu_3295_p2;
    wire   [0:0] icmp_ln133_30_fu_3289_p2;
    wire   [0:0] or_ln133_14_fu_3283_p2;
    wire   [0:0] or_ln133_15_fu_3301_p2;
    wire   [0:0] and_ln133_14_fu_3307_p2;
    wire   [0:0] and_ln133_15_fu_3313_p2;
    wire   [63:0] bitcast_ln134_6_fu_3326_p1;
    wire   [10:0] tmp_71_fu_3329_p4;
    wire   [51:0] trunc_ln134_6_fu_3339_p1;
    wire   [0:0] icmp_ln134_13_fu_3349_p2;
    wire   [0:0] icmp_ln134_12_fu_3343_p2;
    wire   [0:0] or_ln134_6_fu_3355_p2;
    wire   [0:0] and_ln134_13_fu_3361_p2;
    wire   [0:0] and_ln134_14_fu_3367_p2;
    wire   [63:0] bitcast_ln135_14_fu_3380_p1;
    wire   [63:0] bitcast_ln135_15_fu_3397_p1;
    wire   [10:0] tmp_73_fu_3383_p4;
    wire   [51:0] trunc_ln135_14_fu_3393_p1;
    wire   [0:0] icmp_ln135_29_fu_3420_p2;
    wire   [0:0] icmp_ln135_28_fu_3414_p2;
    wire   [10:0] tmp_74_fu_3400_p4;
    wire   [51:0] trunc_ln135_15_fu_3410_p1;
    wire   [0:0] icmp_ln135_31_fu_3438_p2;
    wire   [0:0] icmp_ln135_30_fu_3432_p2;
    wire   [0:0] or_ln135_14_fu_3426_p2;
    wire   [0:0] or_ln135_15_fu_3444_p2;
    wire   [0:0] and_ln135_14_fu_3450_p2;
    wire   [0:0] and_ln135_15_fu_3456_p2;
    wire   [63:0] bitcast_ln136_6_fu_3468_p1;
    wire   [10:0] tmp_76_fu_3471_p4;
    wire   [51:0] trunc_ln136_6_fu_3481_p1;
    wire   [0:0] icmp_ln136_13_fu_3491_p2;
    wire   [0:0] icmp_ln136_12_fu_3485_p2;
    wire   [0:0] or_ln136_6_fu_3497_p2;
    wire   [0:0] and_ln136_13_fu_3503_p2;
    wire   [0:0] and_ln136_14_fu_3509_p2;
    wire   [63:0] bitcast_ln139_fu_3521_p1;
    wire   [63:0] bitcast_ln139_1_fu_3538_p1;
    wire   [10:0] tmp_78_fu_3524_p4;
    wire   [51:0] trunc_ln139_fu_3534_p1;
    wire   [0:0] icmp_ln139_1_fu_3561_p2;
    wire   [0:0] icmp_ln139_fu_3555_p2;
    wire   [10:0] tmp_79_fu_3541_p4;
    wire   [51:0] trunc_ln139_1_fu_3551_p1;
    wire   [0:0] icmp_ln139_3_fu_3579_p2;
    wire   [0:0] icmp_ln139_2_fu_3573_p2;
    wire   [0:0] or_ln139_fu_3567_p2;
    wire   [0:0] or_ln139_1_fu_3585_p2;
    wire   [63:0] bitcast_ln139_2_fu_3597_p1;
    wire   [10:0] tmp_81_fu_3600_p4;
    wire   [51:0] trunc_ln139_2_fu_3610_p1;
    wire   [0:0] icmp_ln139_5_fu_3620_p2;
    wire   [0:0] icmp_ln139_4_fu_3614_p2;
    wire   [0:0] or_ln139_2_fu_3626_p2;
    wire   [0:0] and_ln139_3_fu_3632_p2;
    wire   [63:0] bitcast_ln140_fu_3643_p1;
    wire   [10:0] tmp_83_fu_3646_p4;
    wire   [51:0] trunc_ln140_fu_3656_p1;
    wire   [0:0] icmp_ln140_1_fu_3666_p2;
    wire   [0:0] icmp_ln140_fu_3660_p2;
    wire   [0:0] or_ln140_1_fu_3672_p2;
    wire   [0:0] and_ln140_1_fu_3678_p2;
    wire   [0:0] and_ln140_4_fu_3695_p2;
    wire   [0:0] and_ln141_fu_3700_p2;
    wire   [0:0] and_ln140_2_fu_3684_p2;
    wire   [0:0] or_ln140_fu_3705_p2;
    wire   [0:0] and_ln142_1_fu_3717_p2;
    wire   [0:0] and_ln142_fu_3722_p2;
    wire   [0:0] and_ln139_2_fu_3732_p2;
    wire   [0:0] and_ln139_fu_3736_p2;
    reg   [4:0] grp_fu_807_opcode;
    wire    ap_block_pp0_stage6_00001;
    wire    ap_block_pp0_stage7_00001;
    wire    ap_block_pp0_stage8_00001;
    wire    ap_block_pp0_stage9_00001;
    wire    ap_block_pp0_stage10_00001;
    wire    ap_block_pp0_stage11_00001;
    wire    ap_block_pp0_stage12_00001;
    wire    ap_block_pp0_stage13_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage5_00001;
    reg   [4:0] grp_fu_811_opcode;
    reg   [4:0] grp_fu_815_opcode;
    reg   [13:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to4;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    reg    ap_idle_pp0_0to3;
    reg    ap_reset_idle_pp0;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_enable_pp0;
    wire   [6:0] mul_ln120_fu_972_p00;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 14'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
    end

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1095 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_771_p0),
        .din1(grp_fu_771_p1),
        .ce(1'b1),
        .dout(grp_fu_771_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1096 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_776_p0),
        .din1(grp_fu_776_p1),
        .ce(1'b1),
        .dout(grp_fu_776_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1097 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_781_p0),
        .din1(grp_fu_781_p1),
        .ce(1'b1),
        .dout(grp_fu_781_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1098 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_786_p0),
        .din1(grp_fu_786_p1),
        .ce(1'b1),
        .dout(grp_fu_786_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1099 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_791_p0),
        .din1(grp_fu_791_p1),
        .ce(1'b1),
        .dout(grp_fu_791_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1100 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_795_p0),
        .din1(grp_fu_795_p1),
        .ce(1'b1),
        .dout(grp_fu_795_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1101 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_799_p0),
        .din1(grp_fu_799_p1),
        .ce(1'b1),
        .dout(grp_fu_799_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1102 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_803_p0),
        .din1(grp_fu_803_p1),
        .ce(1'b1),
        .dout(grp_fu_803_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1103 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_807_p0),
        .din1(grp_fu_807_p1),
        .ce(1'b1),
        .opcode(grp_fu_807_opcode),
        .dout(grp_fu_807_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1104 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_811_p0),
        .din1(grp_fu_811_p1),
        .ce(1'b1),
        .opcode(grp_fu_811_opcode),
        .dout(grp_fu_811_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1105 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_815_p0),
        .din1(grp_fu_815_p1),
        .ce(1'b1),
        .opcode(grp_fu_815_opcode),
        .dout(grp_fu_815_p2)
    );

    main_mul_2ns_6ns_7_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(2),
        .din1_WIDTH(6),
        .dout_WIDTH(7)
    ) mul_2ns_6ns_7_1_1_U1106 (
        .din0(mul_ln120_fu_972_p0),
        .din1(mul_ln120_fu_972_p1),
        .dout(mul_ln120_fu_972_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                ap_enable_reg_pp0_iter4 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                reg_835 <= p1_q0;
            end else if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                reg_835 <= p1_q1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13_11001) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                reg_842 <= p1_q0;
            end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                reg_842 <= p1_q1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            reg_849 <= p1_q0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            reg_849 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            add_ln120_2_reg_3786 <= add_ln120_2_fu_1005_p2;
            min2_5_reg_4871 <= min2_5_fu_2369_p3;
            mul_ln120_reg_3751 <= mul_ln120_fu_972_p2;
            p2_offset_cast_reg_3746[2 : 0] <= p2_offset_cast_fu_934_p1[2 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            and_ln135_reg_4740 <= and_ln135_fu_1485_p2;
            max1_reg_4726 <= max1_fu_1391_p3;
            min1_2_reg_4733 <= min1_2_fu_1405_p3;
            mul20_6_2_reg_4626_pp0_iter2_reg <= mul20_6_2_reg_4626;
            mul25_6_2_reg_4631_pp0_iter2_reg <= mul25_6_2_reg_4631;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            and_ln139_1_reg_5036 <= and_ln139_1_fu_3591_p2;
            and_ln139_4_reg_5041 <= and_ln139_4_fu_3638_p2;
            and_ln140_3_reg_5047 <= and_ln140_3_fu_3689_p2;
            and_ln140_reg_5052 <= and_ln140_fu_3711_p2;
            max1_7_reg_4878 <= max1_7_fu_2458_p3;
            max2_7_reg_4897 <= max2_7_fu_2602_p3;
            min1_6_reg_4885 <= min1_6_fu_2512_p3;
            or_ln135_8_reg_4892 <= or_ln135_8_fu_2566_p2;
            p2_0_0_load_reg_3952 <= p2_0_0_q0;
            p2_0_1_load_reg_3957 <= p2_0_1_q0;
            p2_0_2_load_reg_3962 <= p2_0_2_q0;
            p2_1_0_load_reg_3967 <= p2_1_0_q0;
            p2_1_1_load_reg_3972 <= p2_1_1_q0;
            p2_1_2_load_reg_3977 <= p2_1_2_q0;
            p2_2_0_load_reg_3982 <= p2_2_0_q0;
            p2_2_1_load_reg_3987 <= p2_2_1_q0;
            p2_2_2_load_reg_3992 <= p2_2_2_q0;
            p2_3_0_load_reg_3997 <= p2_3_0_q0;
            p2_3_1_load_reg_4002 <= p2_3_1_q0;
            p2_3_2_load_reg_4007 <= p2_3_2_q0;
            p2_4_0_load_reg_4012 <= p2_4_0_q0;
            p2_4_1_load_reg_4017 <= p2_4_1_q0;
            p2_4_2_load_reg_4022 <= p2_4_2_q0;
            p2_5_0_load_reg_4027 <= p2_5_0_q0;
            p2_5_1_load_reg_4032 <= p2_5_1_q0;
            p2_5_2_load_reg_4037 <= p2_5_2_q0;
            p2_6_0_load_reg_4042 <= p2_6_0_q0;
            p2_6_1_load_reg_4047 <= p2_6_1_q0;
            p2_6_2_load_reg_4052 <= p2_6_2_q0;
            p2_7_0_load_reg_4057 <= p2_7_0_q0;
            p2_7_1_load_reg_4062 <= p2_7_1_q0;
            p2_7_2_load_reg_4067 <= p2_7_2_q0;
            p2_8_0_load_reg_4072 <= p2_8_0_q0;
            p2_8_1_load_reg_4077 <= p2_8_1_q0;
            p2_8_2_load_reg_4446 <= p2_8_2_q0;
            sub_ln120_1_reg_3932 <= sub_ln120_1_fu_1036_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            axis_load_1_reg_4105 <= axis_q0;
            axis_load_reg_4097   <= axis_q1;
            p1_load_6_reg_4113   <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            axis_load_2_reg_4128 <= axis_q0;
            p1_load_12_reg_4136  <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            max1_10_reg_4986 <= max1_10_fu_3319_p3;
            max2_reg_4751 <= max2_fu_1495_p3;
            min1_9_reg_4993 <= min1_9_fu_3373_p3;
            min2_2_reg_4758 <= min2_2_fu_1509_p3;
            mul20_7_2_reg_4636_pp0_iter2_reg <= mul20_7_2_reg_4636;
            mul25_7_2_reg_4641_pp0_iter2_reg <= mul25_7_2_reg_4641;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            max1_11_reg_4451 <= grp_fu_771_p2;
            max2_11_reg_4456 <= grp_fu_776_p2;
            mul20_7_reg_4471 <= grp_fu_799_p2;
            mul20_8_reg_4461 <= grp_fu_791_p2;
            mul25_7_reg_4476 <= grp_fu_803_p2;
            mul25_8_reg_4466 <= grp_fu_795_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            max1_1_reg_4646 <= grp_fu_771_p2;
            max2_1_reg_4651 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            max1_4_reg_4779 <= max1_4_fu_1600_p3;
            max2_4_reg_4798 <= max2_4_fu_1744_p3;
            min1_3_reg_4786 <= min1_3_fu_1654_p3;
            or_ln135_2_reg_4793 <= or_ln135_2_fu_1708_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            max1_5_reg_4812 <= max1_5_fu_1887_p3;
            max2_5_reg_4831 <= max2_5_fu_2031_p3;
            min1_4_reg_4819 <= min1_4_fu_1941_p3;
            or_ln135_4_reg_4826 <= or_ln135_4_fu_1995_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            max1_6_reg_4845 <= max1_6_fu_2174_p3;
            max2_6_reg_4864 <= max2_6_fu_2317_p3;
            min1_5_reg_4852 <= min1_5_fu_2228_p3;
            or_ln135_6_reg_4859 <= or_ln135_6_fu_2281_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            max1_8_reg_4920 <= max1_8_fu_2745_p3;
            max2_8_reg_4939 <= max2_8_fu_2889_p3;
            min1_7_reg_4927 <= min1_7_fu_2799_p3;
            or_ln135_10_reg_4934 <= or_ln135_10_fu_2853_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            max1_9_reg_4953 <= max1_9_fu_3032_p3;
            max2_9_reg_4972 <= max2_9_fu_3176_p3;
            min1_8_reg_4960 <= min1_8_fu_3086_p3;
            or_ln135_12_reg_4967 <= or_ln135_12_fu_3140_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            max2_10_reg_5001 <= max2_10_fu_3462_p3;
            min2_3_reg_4805  <= min2_3_fu_1797_p3;
            min2_9_reg_5009  <= min2_9_fu_3515_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            min2_4_reg_4838 <= min2_4_fu_2084_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            min2_6_reg_4913 <= min2_6_fu_2655_p3;
            or_ln140_2_reg_5062 <= or_ln140_2_fu_3727_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            min2_7_reg_4946 <= min2_7_fu_2942_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            min2_8_reg_4979 <= min2_8_fu_3229_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            mul1_reg_4241 <= grp_fu_799_p2;
            mul2_reg_4246 <= grp_fu_803_p2;
            mul6_reg_4236 <= grp_fu_795_p2;
            mul_reg_4231 <= grp_fu_791_p2;
            p1_load_16_reg_4251 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            mul20_1_1_reg_4371 <= grp_fu_791_p2;
            mul20_5_reg_4381 <= grp_fu_799_p2;
            mul25_1_1_reg_4376 <= grp_fu_795_p2;
            mul25_5_reg_4386 <= grp_fu_803_p2;
            p1_load_20_reg_4391 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            mul20_1_2_reg_4491 <= grp_fu_791_p2;
            mul20_4_1_reg_4506 <= grp_fu_799_p2;
            mul25_1_2_reg_4496 <= grp_fu_795_p2;
            mul25_4_1_reg_4511 <= grp_fu_803_p2;
            n1_3_reg_4481 <= grp_fu_771_p2;
            n2_3_reg_4486 <= grp_fu_776_p2;
            n2_6_reg_4501 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            mul20_1_reg_4266 <= grp_fu_791_p2;
            mul20_2_reg_4276 <= grp_fu_799_p2;
            mul25_1_reg_4271 <= grp_fu_795_p2;
            mul25_2_reg_4281 <= grp_fu_803_p2;
            p1_load_19_reg_4286 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            mul20_2_1_reg_4396 <= grp_fu_791_p2;
            mul20_6_reg_4406 <= grp_fu_799_p2;
            mul25_2_1_reg_4401 <= grp_fu_795_p2;
            mul25_6_reg_4411 <= grp_fu_803_p2;
            p1_load_26_reg_4416 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul20_2_2_reg_4516 <= grp_fu_791_p2;
            mul20_5_1_reg_4536 <= grp_fu_799_p2;
            mul25_2_2_reg_4521 <= grp_fu_795_p2;
            mul25_5_1_reg_4541 <= grp_fu_803_p2;
            n1_9_reg_4526 <= grp_fu_771_p2;
            n2_9_reg_4531 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            mul20_3_1_reg_4436 <= grp_fu_799_p2;
            mul25_3_1_reg_4441 <= grp_fu_803_p2;
            mul6_2_reg_4431 <= grp_fu_795_p2;
            mul_2_reg_4426 <= grp_fu_791_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            mul20_3_2_reg_4546 <= grp_fu_791_p2;
            mul20_6_1_reg_4566 <= grp_fu_799_p2;
            mul25_3_2_reg_4551 <= grp_fu_795_p2;
            mul25_6_1_reg_4571 <= grp_fu_803_p2;
            n1_12_reg_4556 <= grp_fu_771_p2;
            n2_12_reg_4561 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            mul20_3_reg_4311 <= grp_fu_799_p2;
            mul25_3_reg_4316 <= grp_fu_803_p2;
            mul6_1_reg_4306 <= grp_fu_795_p2;
            mul_1_reg_4301 <= grp_fu_791_p2;
            p1_load_22_reg_4321 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            mul20_4_2_reg_4576 <= grp_fu_791_p2;
            mul20_7_1_reg_4596 <= grp_fu_799_p2;
            mul25_4_2_reg_4581 <= grp_fu_795_p2;
            mul25_7_1_reg_4601 <= grp_fu_803_p2;
            n1_15_reg_4586 <= grp_fu_771_p2;
            n2_15_reg_4591 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            mul20_4_reg_4346 <= grp_fu_799_p2;
            mul20_s_reg_4336 <= grp_fu_791_p2;
            mul25_4_reg_4351 <= grp_fu_803_p2;
            mul25_s_reg_4341 <= grp_fu_795_p2;
            p1_load_25_reg_4356 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            mul20_5_2_reg_4606 <= grp_fu_791_p2;
            mul20_6_2_reg_4626 <= grp_fu_799_p2;
            mul25_5_2_reg_4611 <= grp_fu_795_p2;
            mul25_6_2_reg_4631 <= grp_fu_803_p2;
            n1_18_reg_4616 <= grp_fu_771_p2;
            n2_18_reg_4621 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            mul20_7_2_reg_4636 <= grp_fu_791_p2;
            mul25_7_2_reg_4641 <= grp_fu_795_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            n1_10_reg_4676 <= grp_fu_771_p2;
            n1_21_reg_4686 <= grp_fu_781_p2;
            n2_10_reg_4681 <= grp_fu_776_p2;
            n2_21_reg_4691 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            n1_13_reg_4696 <= grp_fu_771_p2;
            n2_13_reg_4701 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            n1_16_reg_4706 <= grp_fu_771_p2;
            n2_16_reg_4711 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            n1_19_reg_4716 <= grp_fu_771_p2;
            n2_19_reg_4721 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            n1_22_reg_4774 <= grp_fu_781_p2;
            n2_11_reg_4765 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            n1_4_reg_4656 <= grp_fu_771_p2;
            n1_7_reg_4666 <= grp_fu_781_p2;
            n2_4_reg_4661 <= grp_fu_776_p2;
            n2_7_reg_4671 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            n2_23_reg_4904 <= grp_fu_776_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            p1_load_10_reg_4181 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            p1_load_13_reg_4196 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            p1_load_2_reg_4211 <= p1_q0;
            p1_load_5_reg_4216 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            p1_load_4_reg_4151 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            p1_load_7_reg_4166 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            p1_load_reg_3947 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            reg_819 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_824 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_830 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            reg_855 <= grp_fu_781_p2;
            reg_862 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_869 <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)))) begin
            reg_876 <= grp_fu_781_p2;
            reg_883 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_890 <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_898 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_905 <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_911 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_917 <= grp_fu_786_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_923 <= grp_fu_771_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            tmp_80_reg_5057 <= grp_fu_811_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            tmp_82_reg_5016 <= grp_fu_811_p2;
            tmp_84_reg_5021 <= grp_fu_815_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            tmp_85_reg_5026 <= grp_fu_811_p2;
            tmp_86_reg_5031 <= grp_fu_815_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            tmp_9_reg_4746 <= grp_fu_815_p2;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to3 = 1'b1;
        end else begin
            ap_idle_pp0_0to3 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to4 = 1'b1;
        end else begin
            ap_idle_pp0_1to4 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0_0to3 == 1'b1) & (ap_start == 1'b0))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                axis_address0 = zext_ln120_8_fu_1082_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                axis_address0 = zext_ln120_7_fu_1052_p1;
            end else begin
                axis_address0 = 'bx;
            end
        end else begin
            axis_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            axis_ce0 = 1'b1;
        end else begin
            axis_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            axis_ce1 = 1'b1;
        end else begin
            axis_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_771_p0 = n1_22_reg_4774;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_771_p0 = n1_10_reg_4676;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_771_p0 = n1_18_reg_4616;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_771_p0 = n1_15_reg_4586;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_771_p0 = n1_12_reg_4556;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_771_p0 = n1_9_reg_4526;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_771_p0 = n1_3_reg_4481;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_771_p0 = max1_11_reg_4451;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_771_p0 = mul20_6_reg_4406;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_771_p0 = mul20_5_reg_4381;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_771_p0 = mul20_4_reg_4346;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_771_p0 = mul20_3_reg_4311;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_771_p0 = mul20_1_reg_4266;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_771_p0 = mul_reg_4231;
        end else begin
            grp_fu_771_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_771_p1 = mul20_7_2_reg_4636_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_771_p1 = mul20_3_2_reg_4546;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_771_p1 = mul20_6_1_reg_4566;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_771_p1 = mul20_5_1_reg_4536;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_771_p1 = mul20_4_1_reg_4506;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_771_p1 = mul20_3_1_reg_4436;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_771_p1 = mul20_1_1_reg_4371;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_771_p1 = mul_1_reg_4301;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_771_p1 = 64'd0;
        end else begin
            grp_fu_771_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_776_p0 = reg_898;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_776_p0 = n2_10_reg_4681;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_776_p0 = n2_18_reg_4621;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_776_p0 = n2_15_reg_4591;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_776_p0 = n2_12_reg_4561;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_776_p0 = n2_9_reg_4531;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_776_p0 = n2_3_reg_4486;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_776_p0 = max2_11_reg_4456;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_776_p0 = mul25_6_reg_4411;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_776_p0 = mul25_5_reg_4386;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_776_p0 = mul25_4_reg_4351;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_776_p0 = mul25_3_reg_4316;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_776_p0 = mul25_1_reg_4271;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_776_p0 = mul6_reg_4236;
        end else begin
            grp_fu_776_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_776_p1 = mul25_7_2_reg_4641_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_776_p1 = mul25_3_2_reg_4551;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_776_p1 = mul25_6_1_reg_4571;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_776_p1 = mul25_5_1_reg_4541;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_776_p1 = mul25_4_1_reg_4511;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_776_p1 = mul25_3_1_reg_4441;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_776_p1 = mul25_1_1_reg_4376;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_776_p1 = mul6_1_reg_4306;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_776_p1 = 64'd0;
        end else begin
            grp_fu_776_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_781_p0 = n1_19_reg_4716;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_781_p0 = n1_16_reg_4706;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_781_p0 = n1_13_reg_4696;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_781_p0 = n1_21_reg_4686;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_781_p0 = n1_7_reg_4666;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_781_p0 = n1_4_reg_4656;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_781_p0 = reg_876;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_781_p0 = max1_1_reg_4646;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_781_p0 = mul20_7_reg_4471;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_781_p0 = reg_869;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_781_p0 = reg_855;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_781_p0 = mul20_2_reg_4276;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_781_p0 = mul1_reg_4241;
        end else begin
            grp_fu_781_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_781_p1 = mul20_6_2_reg_4626_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_781_p1 = mul20_5_2_reg_4606;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_781_p1 = mul20_4_2_reg_4576;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_781_p1 = mul20_7_1_reg_4596;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_781_p1 = mul20_2_2_reg_4516;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_781_p1 = mul20_1_2_reg_4491;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_781_p1 = mul20_8_reg_4461;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_781_p1 = mul_2_reg_4426;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_781_p1 = mul20_2_1_reg_4396;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_781_p1 = mul20_s_reg_4336;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_781_p1 = 64'd0;
        end else begin
            grp_fu_781_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_786_p0 = n2_19_reg_4721;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_786_p0 = n2_16_reg_4711;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_786_p0 = n2_13_reg_4701;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_786_p0 = n2_21_reg_4691;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_786_p0 = n2_7_reg_4671;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_786_p0 = n2_4_reg_4661;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_786_p0 = reg_883;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_786_p0 = max2_1_reg_4651;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_786_p0 = mul25_7_reg_4476;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_786_p0 = n2_6_reg_4501;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_786_p0 = reg_862;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_786_p0 = mul25_2_reg_4281;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_786_p0 = mul2_reg_4246;
        end else begin
            grp_fu_786_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_786_p1 = mul25_6_2_reg_4631_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_786_p1 = mul25_5_2_reg_4611;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_786_p1 = mul25_4_2_reg_4581;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_786_p1 = mul25_7_1_reg_4601;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_786_p1 = mul25_2_2_reg_4521;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_786_p1 = mul25_1_2_reg_4496;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_786_p1 = mul25_8_reg_4466;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_786_p1 = mul6_2_reg_4431;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_786_p1 = mul25_2_1_reg_4401;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_786_p1 = mul25_s_reg_4341;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_786_p1 = 64'd0;
        end else begin
            grp_fu_786_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_791_p0 = p1_load_26_reg_4416;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_791_p0 = p1_load_20_reg_4391;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_791_p0 = reg_842;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_791_p0 = reg_835;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_791_p0 = reg_824;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_791_p0 = p1_load_5_reg_4216;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_791_p0 = p1_load_2_reg_4211;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_791_p0 = p1_load_10_reg_4181;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_791_p0 = p1_load_7_reg_4166;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_791_p0 = p1_load_4_reg_4151;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_791_p0 = reg_830;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_791_p0 = p1_load_6_reg_4113;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_791_p0 = p1_load_reg_3947;
        end else begin
            grp_fu_791_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_791_p1 = axis_load_2_reg_4128;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_791_p1 = axis_load_1_reg_4105;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_791_p1 = axis_load_reg_4097;
        end else begin
            grp_fu_791_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_795_p0 = p2_8_2_load_reg_4446;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_795_p0 = p2_6_2_load_reg_4052;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_795_p0 = p2_5_2_load_reg_4037;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_795_p0 = p2_4_2_load_reg_4022;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_795_p0 = p2_3_2_load_reg_4007;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_795_p0 = p2_2_2_load_reg_3992;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_795_p0 = p2_1_2_load_reg_3977;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_795_p0 = p2_0_2_load_reg_3962;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_795_p0 = p2_3_1_load_reg_4002;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_795_p0 = p2_2_1_load_reg_3987;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_795_p0 = p2_1_1_load_reg_3972;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_795_p0 = p2_0_1_load_reg_3957;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_795_p0 = p2_2_0_load_reg_3982;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_795_p0 = p2_0_0_load_reg_3952;
        end else begin
            grp_fu_795_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_795_p1 = axis_load_2_reg_4128;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_795_p1 = axis_load_1_reg_4105;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_795_p1 = axis_load_reg_4097;
        end else begin
            grp_fu_795_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_799_p0 = p1_load_25_reg_4356;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_799_p0 = p1_load_22_reg_4321;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_799_p0 = p1_load_19_reg_4286;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_799_p0 = p1_load_16_reg_4251;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_799_p0 = p1_load_13_reg_4196;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_799_p0 = reg_849;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_799_p0 = reg_842;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_799_p0 = reg_835;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_799_p0 = p1_load_12_reg_4136;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_799_p0 = reg_824;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_799_p0 = reg_819;
        end else begin
            grp_fu_799_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_799_p1 = axis_load_2_reg_4128;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_799_p1 = axis_load_1_reg_4105;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_799_p1 = axis_load_reg_4097;
        end else begin
            grp_fu_799_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_803_p0 = p2_7_2_load_reg_4067;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_803_p0 = p2_8_1_load_reg_4077;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_803_p0 = p2_7_1_load_reg_4062;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_803_p0 = p2_6_1_load_reg_4047;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_803_p0 = p2_5_1_load_reg_4032;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_803_p0 = p2_8_0_load_reg_4072;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_803_p0 = p2_4_1_load_reg_4017;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_803_p0 = p2_7_0_load_reg_4057;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_803_p0 = p2_6_0_load_reg_4042;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_803_p0 = p2_5_0_load_reg_4027;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_803_p0 = p2_4_0_load_reg_4012;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_803_p0 = p2_3_0_load_reg_3997;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_803_p0 = p2_1_0_load_reg_3967;
        end else begin
            grp_fu_803_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_803_p1 = axis_load_2_reg_4128;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_803_p1 = axis_load_1_reg_4105;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_803_p1 = axis_load_reg_4097;
        end else begin
            grp_fu_803_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_807_opcode = 5'd4;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_807_opcode = 5'd2;
        end else begin
            grp_fu_807_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_807_p0 = reg_869;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_807_p0 = reg_862;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_807_p0 = reg_855;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_807_p0 = n2_11_reg_4765;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_807_p0 = reg_923;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_807_p0 = reg_917;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_807_p0 = reg_890;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_807_p0 = reg_911;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_807_p0 = reg_905;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_807_p0 = reg_883;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_807_p0 = reg_876;
        end else begin
            grp_fu_807_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_807_p1 = min2_7_reg_4946;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_807_p1 = max1_8_reg_4920;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_807_p1 = min2_6_reg_4913;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_807_p1 = max1_7_reg_4878;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_807_p1 = min2_5_reg_4871;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_807_p1 = max1_6_reg_4845;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_807_p1 = min2_4_reg_4838;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_807_p1 = max1_5_reg_4812;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_807_p1 = min2_3_reg_4805;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_807_p1 = max1_4_reg_4779;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_807_p1 = min2_2_reg_4758;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_807_p1 = max1_reg_4726;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_807_p1 = reg_898;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_807_p1 = reg_890;
        end else begin
            grp_fu_807_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_811_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_811_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_811_opcode = 5'd2;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_811_opcode = 5'd4;
        end else begin
            grp_fu_811_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_811_p0 = min1_9_reg_4993;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_811_p0 = max1_10_reg_4986;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_811_p0 = n2_23_reg_4904;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_811_p0 = reg_869;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_811_p0 = reg_855;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_811_p0 = reg_923;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_811_p0 = reg_890;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_811_p0 = reg_905;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_811_p0 = reg_876;
        end else begin
            grp_fu_811_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_811_p1 = max2_10_reg_5001;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_811_p1 = min2_9_reg_5009;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_811_p1 = max2_9_reg_4972;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_811_p1 = max1_9_reg_4953;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_811_p1 = min1_7_reg_4927;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_811_p1 = min1_6_reg_4885;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_811_p1 = min1_5_reg_4852;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_811_p1 = min1_4_reg_4819;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_811_p1 = min1_3_reg_4786;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_811_p1 = min1_2_reg_4733;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_811_p1 = reg_890;
        end else begin
            grp_fu_811_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_815_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_815_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_815_opcode = 5'd4;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_815_opcode = 5'd2;
        end else begin
            grp_fu_815_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_815_p0 = min2_9_reg_5009;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_815_p0 = max2_10_reg_5001;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_815_p0 = min1_9_reg_4993;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_815_p0 = n2_23_reg_4904;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_815_p0 = reg_923;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_815_p0 = reg_862;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_815_p0 = n2_11_reg_4765;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_815_p0 = reg_917;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_815_p0 = reg_911;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_815_p0 = reg_883;
        end else begin
            grp_fu_815_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_815_p1 = min1_9_reg_4993;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_815_p1 = max1_10_reg_4986;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_815_p1 = max2_10_reg_5001;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_815_p1 = min2_8_reg_4979;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_815_p1 = min1_8_reg_4960;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_815_p1 = max2_8_reg_4939;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_815_p1 = max2_7_reg_4897;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_815_p1 = max2_6_reg_4864;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_815_p1 = max2_5_reg_4831;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_815_p1 = max2_4_reg_4798;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_815_p1 = max2_fu_1495_p3;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_815_p1 = reg_898;
        end else begin
            grp_fu_815_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address0 = zext_ln129_20_fu_1292_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address0 = zext_ln129_14_fu_1272_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address0 = zext_ln129_11_fu_1252_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address0 = zext_ln129_8_fu_1232_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address0 = zext_ln129_5_fu_1212_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address0 = zext_ln129_13_fu_1192_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address0 = zext_ln120_4_fu_1172_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address0 = zext_ln129_10_fu_1152_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address0 = zext_ln129_7_fu_1132_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address0 = zext_ln129_4_fu_1112_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address0 = zext_ln120_3_fu_1092_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address0 = zext_ln129_6_fu_1062_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address0 = zext_ln129_3_fu_1026_p1;
            end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                p1_address0 = zext_ln120_2_fu_978_p1;
            end else begin
                p1_address0 = 'bx;
            end
        end else begin
            p1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address1 = zext_ln129_23_fu_1302_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address1 = zext_ln129_17_fu_1282_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address1 = zext_ln129_22_fu_1262_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address1 = zext_ln129_19_fu_1242_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address1 = zext_ln129_16_fu_1222_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address1 = zext_ln129_21_fu_1202_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address1 = zext_ln129_2_fu_1182_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address1 = zext_ln129_18_fu_1162_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address1 = zext_ln129_15_fu_1142_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address1 = zext_ln129_12_fu_1122_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address1 = zext_ln129_1_fu_1102_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address1 = zext_ln129_9_fu_1072_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address1 = zext_ln129_fu_1016_p1;
            end else begin
                p1_address1 = 'bx;
            end
        end else begin
            p1_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            p1_ce0 = 1'b1;
        end else begin
            p1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            p1_ce1 = 1'b1;
        end else begin
            p1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_0_ce0 = 1'b1;
        end else begin
            p2_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_1_ce0 = 1'b1;
        end else begin
            p2_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_2_ce0 = 1'b1;
        end else begin
            p2_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_0_ce0 = 1'b1;
        end else begin
            p2_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_1_ce0 = 1'b1;
        end else begin
            p2_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_2_ce0 = 1'b1;
        end else begin
            p2_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_0_ce0 = 1'b1;
        end else begin
            p2_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_1_ce0 = 1'b1;
        end else begin
            p2_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_2_ce0 = 1'b1;
        end else begin
            p2_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_0_ce0 = 1'b1;
        end else begin
            p2_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_1_ce0 = 1'b1;
        end else begin
            p2_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_2_ce0 = 1'b1;
        end else begin
            p2_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_0_ce0 = 1'b1;
        end else begin
            p2_4_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_1_ce0 = 1'b1;
        end else begin
            p2_4_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_2_ce0 = 1'b1;
        end else begin
            p2_4_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_0_ce0 = 1'b1;
        end else begin
            p2_5_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_1_ce0 = 1'b1;
        end else begin
            p2_5_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_2_ce0 = 1'b1;
        end else begin
            p2_5_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_0_ce0 = 1'b1;
        end else begin
            p2_6_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_1_ce0 = 1'b1;
        end else begin
            p2_6_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_2_ce0 = 1'b1;
        end else begin
            p2_6_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_0_ce0 = 1'b1;
        end else begin
            p2_7_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_1_ce0 = 1'b1;
        end else begin
            p2_7_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_2_ce0 = 1'b1;
        end else begin
            p2_7_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_0_ce0 = 1'b1;
        end else begin
            p2_8_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_1_ce0 = 1'b1;
        end else begin
            p2_8_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_2_ce0 = 1'b1;
        end else begin
            p2_8_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_idle_pp0_1to4 == 1'b1) & (ap_start == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_reset_idle_pp0 == 1'b0))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_reset_idle_pp0 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln120_1_fu_1167_p2 = (mul_ln120_reg_3751 + 7'd2);

    assign add_ln120_2_fu_1005_p2 = ($signed(
        sext_ln120_fu_1001_p1
    ) + $signed(
        axis_offset1_cast4_fu_930_p1
    ));

    assign add_ln120_3_fu_1046_p2 = (sub_ln120_1_fu_1036_p2 + 6'd1);

    assign add_ln120_4_fu_1077_p2 = (sub_ln120_1_reg_3932 + 6'd2);

    assign add_ln120_fu_1087_p2 = (mul_ln120_reg_3751 + 7'd1);

    assign add_ln129_10_fu_1147_p2 = (mul_ln120_reg_3751 + 7'd13);

    assign add_ln129_11_fu_1247_p2 = (mul_ln120_reg_3751 + 7'd14);

    assign add_ln129_12_fu_1117_p2 = (mul_ln120_reg_3751 + 7'd15);

    assign add_ln129_13_fu_1187_p2 = (mul_ln120_reg_3751 + 7'd16);

    assign add_ln129_14_fu_1267_p2 = (mul_ln120_reg_3751 + 7'd17);

    assign add_ln129_15_fu_1137_p2 = (mul_ln120_reg_3751 + 7'd18);

    assign add_ln129_16_fu_1217_p2 = (mul_ln120_reg_3751 + 7'd19);

    assign add_ln129_17_fu_1277_p2 = (mul_ln120_reg_3751 + 7'd20);

    assign add_ln129_18_fu_1157_p2 = (mul_ln120_reg_3751 + 7'd21);

    assign add_ln129_19_fu_1237_p2 = (mul_ln120_reg_3751 + 7'd22);

    assign add_ln129_1_fu_1097_p2 = (mul_ln120_reg_3751 + 7'd4);

    assign add_ln129_20_fu_1287_p2 = (mul_ln120_reg_3751 + 7'd23);

    assign add_ln129_21_fu_1197_p2 = (mul_ln120_reg_3751 + 7'd24);

    assign add_ln129_22_fu_1257_p2 = (mul_ln120_reg_3751 + 7'd25);

    assign add_ln129_23_fu_1297_p2 = (mul_ln120_reg_3751 + 7'd26);

    assign add_ln129_2_fu_1177_p2 = (mul_ln120_reg_3751 + 7'd5);

    assign add_ln129_3_fu_1021_p2 = (mul_ln120_reg_3751 + 7'd6);

    assign add_ln129_4_fu_1107_p2 = (mul_ln120_reg_3751 + 7'd7);

    assign add_ln129_5_fu_1207_p2 = (mul_ln120_reg_3751 + 7'd8);

    assign add_ln129_6_fu_1057_p2 = (mul_ln120_reg_3751 + 7'd9);

    assign add_ln129_7_fu_1127_p2 = (mul_ln120_reg_3751 + 7'd10);

    assign add_ln129_8_fu_1227_p2 = (mul_ln120_reg_3751 + 7'd11);

    assign add_ln129_9_fu_1067_p2 = (mul_ln120_reg_3751 + 7'd12);

    assign add_ln129_fu_1011_p2 = (mul_ln120_reg_3751 + 7'd3);

    assign and_ln133_10_fu_2733_p2 = (or_ln133_11_fu_2727_p2 & or_ln133_10_fu_2709_p2);

    assign and_ln133_11_fu_2739_p2 = (grp_fu_807_p2 & and_ln133_10_fu_2733_p2);

    assign and_ln133_12_fu_3020_p2 = (or_ln133_13_fu_3014_p2 & or_ln133_12_fu_2996_p2);

    assign and_ln133_13_fu_3026_p2 = (grp_fu_807_p2 & and_ln133_12_fu_3020_p2);

    assign and_ln133_14_fu_3307_p2 = (or_ln133_15_fu_3301_p2 & or_ln133_14_fu_3283_p2);

    assign and_ln133_15_fu_3313_p2 = (grp_fu_811_p2 & and_ln133_14_fu_3307_p2);

    assign and_ln133_1_fu_1385_p2 = (grp_fu_807_p2 & and_ln133_fu_1379_p2);

    assign and_ln133_2_fu_1588_p2 = (or_ln133_3_fu_1582_p2 & or_ln133_2_fu_1564_p2);

    assign and_ln133_3_fu_1594_p2 = (grp_fu_807_p2 & and_ln133_2_fu_1588_p2);

    assign and_ln133_4_fu_1875_p2 = (or_ln133_5_fu_1869_p2 & or_ln133_4_fu_1851_p2);

    assign and_ln133_5_fu_1881_p2 = (grp_fu_807_p2 & and_ln133_4_fu_1875_p2);

    assign and_ln133_6_fu_2162_p2 = (or_ln133_7_fu_2156_p2 & or_ln133_6_fu_2138_p2);

    assign and_ln133_7_fu_2168_p2 = (grp_fu_807_p2 & and_ln133_6_fu_2162_p2);

    assign and_ln133_8_fu_2446_p2 = (or_ln133_9_fu_2440_p2 & or_ln133_8_fu_2422_p2);

    assign and_ln133_9_fu_2452_p2 = (grp_fu_807_p2 & and_ln133_8_fu_2446_p2);

    assign and_ln133_fu_1379_p2 = (or_ln133_fu_1355_p2 & or_ln133_1_fu_1373_p2);

    assign and_ln134_10_fu_2793_p2 = (grp_fu_811_p2 & and_ln134_9_fu_2787_p2);

    assign and_ln134_11_fu_3074_p2 = (or_ln134_5_fu_3068_p2 & or_ln133_12_fu_2996_p2);

    assign and_ln134_12_fu_3080_p2 = (grp_fu_811_p2 & and_ln134_11_fu_3074_p2);

    assign and_ln134_13_fu_3361_p2 = (or_ln134_6_fu_3355_p2 & or_ln133_14_fu_3283_p2);

    assign and_ln134_14_fu_3367_p2 = (grp_fu_815_p2 & and_ln134_13_fu_3361_p2);

    assign and_ln134_1_fu_1642_p2 = (or_ln134_fu_1636_p2 & or_ln133_2_fu_1564_p2);

    assign and_ln134_2_fu_1648_p2 = (grp_fu_811_p2 & and_ln134_1_fu_1642_p2);

    assign and_ln134_3_fu_1929_p2 = (or_ln134_1_fu_1923_p2 & or_ln133_4_fu_1851_p2);

    assign and_ln134_4_fu_1935_p2 = (grp_fu_811_p2 & and_ln134_3_fu_1929_p2);

    assign and_ln134_5_fu_2216_p2 = (or_ln134_2_fu_2210_p2 & or_ln133_6_fu_2138_p2);

    assign and_ln134_6_fu_2222_p2 = (grp_fu_811_p2 & and_ln134_5_fu_2216_p2);

    assign and_ln134_7_fu_2500_p2 = (or_ln134_3_fu_2494_p2 & or_ln133_8_fu_2422_p2);

    assign and_ln134_8_fu_2506_p2 = (grp_fu_811_p2 & and_ln134_7_fu_2500_p2);

    assign and_ln134_9_fu_2787_p2 = (or_ln134_4_fu_2781_p2 & or_ln133_10_fu_2709_p2);

    assign and_ln134_fu_1399_p2 = (grp_fu_811_p2 & and_ln133_fu_1379_p2);

    assign and_ln135_10_fu_2877_p2 = (or_ln135_11_fu_2871_p2 & or_ln135_10_fu_2853_p2);

    assign and_ln135_11_fu_2883_p2 = (grp_fu_815_p2 & and_ln135_10_fu_2877_p2);

    assign and_ln135_12_fu_3164_p2 = (or_ln135_13_fu_3158_p2 & or_ln135_12_fu_3140_p2);

    assign and_ln135_13_fu_3170_p2 = (grp_fu_815_p2 & and_ln135_12_fu_3164_p2);

    assign and_ln135_14_fu_3450_p2 = (or_ln135_15_fu_3444_p2 & or_ln135_14_fu_3426_p2);

    assign and_ln135_15_fu_3456_p2 = (grp_fu_811_p2 & and_ln135_14_fu_3450_p2);

    assign and_ln135_1_fu_1491_p2 = (tmp_9_reg_4746 & and_ln135_reg_4740);

    assign and_ln135_2_fu_1732_p2 = (or_ln135_3_fu_1726_p2 & or_ln135_2_fu_1708_p2);

    assign and_ln135_3_fu_1738_p2 = (grp_fu_815_p2 & and_ln135_2_fu_1732_p2);

    assign and_ln135_4_fu_2019_p2 = (or_ln135_5_fu_2013_p2 & or_ln135_4_fu_1995_p2);

    assign and_ln135_5_fu_2025_p2 = (grp_fu_815_p2 & and_ln135_4_fu_2019_p2);

    assign and_ln135_6_fu_2305_p2 = (or_ln135_7_fu_2299_p2 & or_ln135_6_fu_2281_p2);

    assign and_ln135_7_fu_2311_p2 = (grp_fu_815_p2 & and_ln135_6_fu_2305_p2);

    assign and_ln135_8_fu_2590_p2 = (or_ln135_9_fu_2584_p2 & or_ln135_8_fu_2566_p2);

    assign and_ln135_9_fu_2596_p2 = (grp_fu_815_p2 & and_ln135_8_fu_2590_p2);

    assign and_ln135_fu_1485_p2 = (or_ln135_fu_1461_p2 & or_ln135_1_fu_1479_p2);

    assign and_ln136_10_fu_2936_p2 = (grp_fu_807_p2 & and_ln136_9_fu_2931_p2);

    assign and_ln136_11_fu_3218_p2 = (or_ln136_5_fu_3212_p2 & or_ln135_12_reg_4967);

    assign and_ln136_12_fu_3223_p2 = (grp_fu_807_p2 & and_ln136_11_fu_3218_p2);

    assign and_ln136_13_fu_3503_p2 = (or_ln136_6_fu_3497_p2 & or_ln135_14_fu_3426_p2);

    assign and_ln136_14_fu_3509_p2 = (grp_fu_815_p2 & and_ln136_13_fu_3503_p2);

    assign and_ln136_1_fu_1786_p2 = (or_ln136_fu_1780_p2 & or_ln135_2_reg_4793);

    assign and_ln136_2_fu_1791_p2 = (grp_fu_807_p2 & and_ln136_1_fu_1786_p2);

    assign and_ln136_3_fu_2073_p2 = (or_ln136_1_fu_2067_p2 & or_ln135_4_reg_4826);

    assign and_ln136_4_fu_2078_p2 = (grp_fu_807_p2 & and_ln136_3_fu_2073_p2);

    assign and_ln136_5_fu_2358_p2 = (or_ln136_2_fu_2352_p2 & or_ln135_6_reg_4859);

    assign and_ln136_6_fu_2363_p2 = (grp_fu_807_p2 & and_ln136_5_fu_2358_p2);

    assign and_ln136_7_fu_2644_p2 = (or_ln136_3_fu_2638_p2 & or_ln135_8_reg_4892);

    assign and_ln136_8_fu_2649_p2 = (grp_fu_807_p2 & and_ln136_7_fu_2644_p2);

    assign and_ln136_9_fu_2931_p2 = (or_ln136_4_fu_2925_p2 & or_ln135_10_reg_4934);

    assign and_ln136_fu_1504_p2 = (grp_fu_807_p2 & and_ln135_reg_4740);

    assign and_ln139_1_fu_3591_p2 = (or_ln139_fu_3567_p2 & or_ln139_1_fu_3585_p2);

    assign and_ln139_2_fu_3732_p2 = (tmp_80_reg_5057 & and_ln139_1_reg_5036);

    assign and_ln139_3_fu_3632_p2 = (or_ln139_fu_3567_p2 & or_ln139_2_fu_3626_p2);

    assign and_ln139_4_fu_3638_p2 = (tmp_82_reg_5016 & and_ln139_3_fu_3632_p2);

    assign and_ln139_fu_3736_p2 = (and_ln139_4_reg_5041 & and_ln139_2_fu_3732_p2);

    assign and_ln140_1_fu_3678_p2 = (or_ln140_1_fu_3672_p2 & or_ln139_1_fu_3585_p2);

    assign and_ln140_2_fu_3684_p2 = (tmp_84_reg_5021 & and_ln140_1_fu_3678_p2);

    assign and_ln140_3_fu_3689_p2 = (or_ln140_1_fu_3672_p2 & or_ln139_2_fu_3626_p2);

    assign and_ln140_4_fu_3695_p2 = (tmp_85_reg_5026 & and_ln140_3_fu_3689_p2);

    assign and_ln140_fu_3711_p2 = (or_ln140_fu_3705_p2 & and_ln140_2_fu_3684_p2);

    assign and_ln141_fu_3700_p2 = (tmp_86_reg_5031 & and_ln139_1_fu_3591_p2);

    assign and_ln142_1_fu_3717_p2 = (grp_fu_815_p2 & and_ln140_3_reg_5047);

    assign and_ln142_fu_3722_p2 = (and_ln142_1_fu_3717_p2 & and_ln139_4_reg_5041);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_return = (or_ln140_2_reg_5062 | and_ln139_fu_3736_p2);

    assign axis_address1 = zext_ln120_6_fu_1041_p1;

    assign axis_offset1_cast4_fu_930_p1 = axis_offset1;

    assign bitcast_ln133_10_fu_2662_p1 = reg_869;

    assign bitcast_ln133_11_fu_2680_p1 = max1_7_reg_4878;

    assign bitcast_ln133_12_fu_2949_p1 = reg_905;

    assign bitcast_ln133_13_fu_2967_p1 = max1_8_reg_4920;

    assign bitcast_ln133_14_fu_3236_p1 = reg_923;

    assign bitcast_ln133_15_fu_3254_p1 = max1_9_reg_4953;

    assign bitcast_ln133_1_fu_1325_p1 = reg_890;

    assign bitcast_ln133_2_fu_1517_p1 = reg_905;

    assign bitcast_ln133_3_fu_1535_p1 = max1_reg_4726;

    assign bitcast_ln133_4_fu_1804_p1 = reg_890;

    assign bitcast_ln133_5_fu_1822_p1 = max1_4_reg_4779;

    assign bitcast_ln133_6_fu_2091_p1 = reg_923;

    assign bitcast_ln133_7_fu_2109_p1 = max1_5_reg_4812;

    assign bitcast_ln133_8_fu_2375_p1 = reg_855;

    assign bitcast_ln133_9_fu_2393_p1 = max1_6_reg_4845;

    assign bitcast_ln133_fu_1307_p1 = reg_876;

    assign bitcast_ln134_1_fu_1894_p1 = min1_3_reg_4786;

    assign bitcast_ln134_2_fu_2181_p1 = min1_4_reg_4819;

    assign bitcast_ln134_3_fu_2465_p1 = min1_5_reg_4852;

    assign bitcast_ln134_4_fu_2752_p1 = min1_6_reg_4885;

    assign bitcast_ln134_5_fu_3039_p1 = min1_7_reg_4927;

    assign bitcast_ln134_6_fu_3326_p1 = min1_8_reg_4960;

    assign bitcast_ln134_fu_1607_p1 = min1_2_reg_4733;

    assign bitcast_ln135_10_fu_2806_p1 = reg_911;

    assign bitcast_ln135_11_fu_2824_p1 = max2_7_reg_4897;

    assign bitcast_ln135_12_fu_3093_p1 = reg_917;

    assign bitcast_ln135_13_fu_3111_p1 = max2_8_reg_4939;

    assign bitcast_ln135_14_fu_3380_p1 = n2_23_reg_4904;

    assign bitcast_ln135_15_fu_3397_p1 = max2_9_reg_4972;

    assign bitcast_ln135_1_fu_1431_p1 = reg_898;

    assign bitcast_ln135_2_fu_1661_p1 = reg_911;

    assign bitcast_ln135_3_fu_1679_p1 = max2_reg_4751;

    assign bitcast_ln135_4_fu_1948_p1 = reg_917;

    assign bitcast_ln135_5_fu_1966_p1 = max2_4_reg_4798;

    assign bitcast_ln135_6_fu_2235_p1 = n2_11_reg_4765;

    assign bitcast_ln135_7_fu_2252_p1 = max2_5_reg_4831;

    assign bitcast_ln135_8_fu_2519_p1 = reg_862;

    assign bitcast_ln135_9_fu_2537_p1 = max2_6_reg_4864;

    assign bitcast_ln135_fu_1413_p1 = reg_883;

    assign bitcast_ln136_1_fu_2038_p1 = min2_3_reg_4805;

    assign bitcast_ln136_2_fu_2323_p1 = min2_4_reg_4838;

    assign bitcast_ln136_3_fu_2609_p1 = min2_5_reg_4871;

    assign bitcast_ln136_4_fu_2896_p1 = min2_6_reg_4913;

    assign bitcast_ln136_5_fu_3183_p1 = min2_7_reg_4946;

    assign bitcast_ln136_6_fu_3468_p1 = min2_8_reg_4979;

    assign bitcast_ln136_fu_1751_p1 = min2_2_reg_4758;

    assign bitcast_ln139_1_fu_3538_p1 = max2_10_reg_5001;

    assign bitcast_ln139_2_fu_3597_p1 = min2_9_reg_5009;

    assign bitcast_ln139_fu_3521_p1 = max1_10_reg_4986;

    assign bitcast_ln140_fu_3643_p1 = min1_9_reg_4993;

    assign icmp_ln133_10_fu_1857_p2 = ((tmp_19_fu_1825_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_11_fu_1863_p2 = ((trunc_ln133_5_fu_1835_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_12_fu_2126_p2 = ((tmp_28_fu_2095_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_13_fu_2132_p2 = ((trunc_ln133_6_fu_2105_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_14_fu_2144_p2 = ((tmp_29_fu_2112_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_15_fu_2150_p2 = ((trunc_ln133_7_fu_2122_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_16_fu_2410_p2 = ((tmp_38_fu_2379_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_17_fu_2416_p2 = ((trunc_ln133_8_fu_2389_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_18_fu_2428_p2 = ((tmp_39_fu_2396_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_19_fu_2434_p2 = ((trunc_ln133_9_fu_2406_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_1_fu_1349_p2 = ((trunc_ln133_fu_1321_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_20_fu_2697_p2 = ((tmp_48_fu_2666_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_21_fu_2703_p2 = ((trunc_ln133_10_fu_2676_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_22_fu_2715_p2 = ((tmp_49_fu_2683_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_23_fu_2721_p2 = ((trunc_ln133_11_fu_2693_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_24_fu_2984_p2 = ((tmp_58_fu_2953_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_25_fu_2990_p2 = ((trunc_ln133_12_fu_2963_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_26_fu_3002_p2 = ((tmp_59_fu_2970_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_27_fu_3008_p2 = ((trunc_ln133_13_fu_2980_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_28_fu_3271_p2 = ((tmp_68_fu_3240_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_29_fu_3277_p2 = ((trunc_ln133_14_fu_3250_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_2_fu_1361_p2 = ((tmp_2_fu_1329_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_30_fu_3289_p2 = ((tmp_69_fu_3257_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_31_fu_3295_p2 = ((trunc_ln133_15_fu_3267_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_3_fu_1367_p2 = ((trunc_ln133_1_fu_1339_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_4_fu_1552_p2 = ((tmp_4_fu_1521_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_5_fu_1558_p2 = ((trunc_ln133_2_fu_1531_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_6_fu_1570_p2 = ((tmp_5_fu_1538_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_7_fu_1576_p2 = ((trunc_ln133_3_fu_1548_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_8_fu_1839_p2 = ((tmp_18_fu_1808_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_9_fu_1845_p2 = ((trunc_ln133_4_fu_1818_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_fu_1343_p2 = ((tmp_1_fu_1311_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_10_fu_3056_p2 = ((tmp_61_fu_3042_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_11_fu_3062_p2 = ((trunc_ln134_5_fu_3052_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_12_fu_3343_p2 = ((tmp_71_fu_3329_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_13_fu_3349_p2 = ((trunc_ln134_6_fu_3339_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_1_fu_1630_p2 = ((trunc_ln134_fu_1620_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_2_fu_1911_p2 = ((tmp_21_fu_1897_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_3_fu_1917_p2 = ((trunc_ln134_1_fu_1907_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_4_fu_2198_p2 = ((tmp_31_fu_2184_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_5_fu_2204_p2 = ((trunc_ln134_2_fu_2194_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_6_fu_2482_p2 = ((tmp_41_fu_2468_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_7_fu_2488_p2 = ((trunc_ln134_3_fu_2478_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_8_fu_2769_p2 = ((tmp_51_fu_2755_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_9_fu_2775_p2 = ((trunc_ln134_4_fu_2765_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_fu_1624_p2 = ((tmp_11_fu_1610_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_10_fu_2001_p2 = ((tmp_24_fu_1969_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_11_fu_2007_p2 = ((trunc_ln135_5_fu_1979_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_12_fu_2269_p2 = ((tmp_33_fu_2238_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_13_fu_2275_p2 = ((trunc_ln135_6_fu_2248_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_14_fu_2287_p2 = ((tmp_34_fu_2255_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_15_fu_2293_p2 = ((trunc_ln135_7_fu_2265_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_16_fu_2554_p2 = ((tmp_43_fu_2523_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_17_fu_2560_p2 = ((trunc_ln135_8_fu_2533_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_18_fu_2572_p2 = ((tmp_44_fu_2540_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_19_fu_2578_p2 = ((trunc_ln135_9_fu_2550_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_1_fu_1455_p2 = ((trunc_ln135_fu_1427_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_20_fu_2841_p2 = ((tmp_53_fu_2810_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_21_fu_2847_p2 = ((trunc_ln135_10_fu_2820_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_22_fu_2859_p2 = ((tmp_54_fu_2827_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_23_fu_2865_p2 = ((trunc_ln135_11_fu_2837_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_24_fu_3128_p2 = ((tmp_63_fu_3097_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_25_fu_3134_p2 = ((trunc_ln135_12_fu_3107_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_26_fu_3146_p2 = ((tmp_64_fu_3114_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_27_fu_3152_p2 = ((trunc_ln135_13_fu_3124_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_28_fu_3414_p2 = ((tmp_73_fu_3383_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_29_fu_3420_p2 = ((trunc_ln135_14_fu_3393_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_2_fu_1467_p2 = ((tmp_8_fu_1435_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_30_fu_3432_p2 = ((tmp_74_fu_3400_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_31_fu_3438_p2 = ((trunc_ln135_15_fu_3410_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_3_fu_1473_p2 = ((trunc_ln135_1_fu_1445_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_4_fu_1696_p2 = ((tmp_13_fu_1665_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_5_fu_1702_p2 = ((trunc_ln135_2_fu_1675_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_6_fu_1714_p2 = ((tmp_14_fu_1682_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_7_fu_1720_p2 = ((trunc_ln135_3_fu_1692_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_8_fu_1983_p2 = ((tmp_23_fu_1952_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_9_fu_1989_p2 = ((trunc_ln135_4_fu_1962_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_fu_1449_p2 = ((tmp_7_fu_1417_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_10_fu_3200_p2 = ((tmp_66_fu_3186_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_11_fu_3206_p2 = ((trunc_ln136_5_fu_3196_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_12_fu_3485_p2 = ((tmp_76_fu_3471_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_13_fu_3491_p2 = ((trunc_ln136_6_fu_3481_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_1_fu_1774_p2 = ((trunc_ln136_fu_1764_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_2_fu_2055_p2 = ((tmp_26_fu_2041_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_3_fu_2061_p2 = ((trunc_ln136_1_fu_2051_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_4_fu_2340_p2 = ((tmp_36_fu_2326_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_5_fu_2346_p2 = ((trunc_ln136_2_fu_2336_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_6_fu_2626_p2 = ((tmp_46_fu_2612_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_7_fu_2632_p2 = ((trunc_ln136_3_fu_2622_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_8_fu_2913_p2 = ((tmp_56_fu_2899_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_9_fu_2919_p2 = ((trunc_ln136_4_fu_2909_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_fu_1768_p2 = ((tmp_16_fu_1754_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_1_fu_3561_p2 = ((trunc_ln139_fu_3534_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_2_fu_3573_p2 = ((tmp_79_fu_3541_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_3_fu_3579_p2 = ((trunc_ln139_1_fu_3551_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_4_fu_3614_p2 = ((tmp_81_fu_3600_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_5_fu_3620_p2 = ((trunc_ln139_2_fu_3610_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_fu_3555_p2 = ((tmp_78_fu_3524_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln140_1_fu_3666_p2 = ((trunc_ln140_fu_3656_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln140_fu_3660_p2 = ((tmp_83_fu_3646_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign max1_10_fu_3319_p3 = ((and_ln133_15_fu_3313_p2[0:0] == 1'b1) ? reg_923 : max1_9_reg_4953);

    assign max1_4_fu_1600_p3 = ((and_ln133_3_fu_1594_p2[0:0] == 1'b1) ? reg_905 : max1_reg_4726);

    assign max1_5_fu_1887_p3 = ((and_ln133_5_fu_1881_p2[0:0] == 1'b1) ? reg_890 : max1_4_reg_4779);

    assign max1_6_fu_2174_p3 = ((and_ln133_7_fu_2168_p2[0:0] == 1'b1) ? reg_923 : max1_5_reg_4812);

    assign max1_7_fu_2458_p3 = ((and_ln133_9_fu_2452_p2[0:0] == 1'b1) ? reg_855 : max1_6_reg_4845);

    assign max1_8_fu_2745_p3 = ((and_ln133_11_fu_2739_p2[0:0] == 1'b1) ? reg_869 : max1_7_reg_4878);

    assign max1_9_fu_3032_p3 = ((and_ln133_13_fu_3026_p2[0:0] == 1'b1) ? reg_905 : max1_8_reg_4920);

    assign max1_fu_1391_p3 = ((and_ln133_1_fu_1385_p2[0:0] == 1'b1) ? reg_876 : reg_890);

    assign max2_10_fu_3462_p3 = ((and_ln135_15_fu_3456_p2[0:0] == 1'b1) ? n2_23_reg_4904 : max2_9_reg_4972);

    assign max2_4_fu_1744_p3 = ((and_ln135_3_fu_1738_p2[0:0] == 1'b1) ? reg_911 : max2_reg_4751);

    assign max2_5_fu_2031_p3 = ((and_ln135_5_fu_2025_p2[0:0] == 1'b1) ? reg_917 : max2_4_reg_4798);

    assign max2_6_fu_2317_p3 = ((and_ln135_7_fu_2311_p2[0:0] == 1'b1) ? n2_11_reg_4765 : max2_5_reg_4831);

    assign max2_7_fu_2602_p3 = ((and_ln135_9_fu_2596_p2[0:0] == 1'b1) ? reg_862 : max2_6_reg_4864);

    assign max2_8_fu_2889_p3 = ((and_ln135_11_fu_2883_p2[0:0] == 1'b1) ? reg_911 : max2_7_reg_4897);

    assign max2_9_fu_3176_p3 = ((and_ln135_13_fu_3170_p2[0:0] == 1'b1) ? reg_917 : max2_8_reg_4939);

    assign max2_fu_1495_p3 = ((and_ln135_1_fu_1491_p2[0:0] == 1'b1) ? reg_883 : reg_898);

    assign min1_2_fu_1405_p3 = ((and_ln134_fu_1399_p2[0:0] == 1'b1) ? reg_876 : reg_890);

    assign min1_3_fu_1654_p3 = ((and_ln134_2_fu_1648_p2[0:0] == 1'b1) ? reg_905 : min1_2_reg_4733);

    assign min1_4_fu_1941_p3 = ((and_ln134_4_fu_1935_p2[0:0] == 1'b1) ? reg_890 : min1_3_reg_4786);

    assign min1_5_fu_2228_p3 = ((and_ln134_6_fu_2222_p2[0:0] == 1'b1) ? reg_923 : min1_4_reg_4819);

    assign min1_6_fu_2512_p3 = ((and_ln134_8_fu_2506_p2[0:0] == 1'b1) ? reg_855 : min1_5_reg_4852);

    assign min1_7_fu_2799_p3 = ((and_ln134_10_fu_2793_p2[0:0] == 1'b1) ? reg_869 : min1_6_reg_4885);

    assign min1_8_fu_3086_p3 = ((and_ln134_12_fu_3080_p2[0:0] == 1'b1) ? reg_905 : min1_7_reg_4927);

    assign min1_9_fu_3373_p3 = ((and_ln134_14_fu_3367_p2[0:0] == 1'b1) ? reg_923 : min1_8_reg_4960);

    assign min2_2_fu_1509_p3 = ((and_ln136_fu_1504_p2[0:0] == 1'b1) ? reg_883 : reg_898);

    assign min2_3_fu_1797_p3 = ((and_ln136_2_fu_1791_p2[0:0] == 1'b1) ? reg_911 : min2_2_reg_4758);

    assign min2_4_fu_2084_p3 = ((and_ln136_4_fu_2078_p2[0:0] == 1'b1) ? reg_917 : min2_3_reg_4805);

    assign min2_5_fu_2369_p3 = ((and_ln136_6_fu_2363_p2[0:0] == 1'b1) ? n2_11_reg_4765 : min2_4_reg_4838);

    assign min2_6_fu_2655_p3 = ((and_ln136_8_fu_2649_p2[0:0] == 1'b1) ? reg_862 : min2_5_reg_4871);

    assign min2_7_fu_2942_p3 = ((and_ln136_10_fu_2936_p2[0:0] == 1'b1) ? reg_911 : min2_6_reg_4913);

    assign min2_8_fu_3229_p3 = ((and_ln136_12_fu_3223_p2[0:0] == 1'b1) ? reg_917 : min2_7_reg_4946);

    assign min2_9_fu_3515_p3 = ((and_ln136_14_fu_3509_p2[0:0] == 1'b1) ? n2_23_reg_4904 : min2_8_reg_4979);

    assign mul_ln120_fu_972_p0 = mul_ln120_fu_972_p00;

    assign mul_ln120_fu_972_p00 = p1_offset;

    assign mul_ln120_fu_972_p1 = 7'd27;

    assign or_ln133_10_fu_2709_p2 = (icmp_ln133_21_fu_2703_p2 | icmp_ln133_20_fu_2697_p2);

    assign or_ln133_11_fu_2727_p2 = (icmp_ln133_23_fu_2721_p2 | icmp_ln133_22_fu_2715_p2);

    assign or_ln133_12_fu_2996_p2 = (icmp_ln133_25_fu_2990_p2 | icmp_ln133_24_fu_2984_p2);

    assign or_ln133_13_fu_3014_p2 = (icmp_ln133_27_fu_3008_p2 | icmp_ln133_26_fu_3002_p2);

    assign or_ln133_14_fu_3283_p2 = (icmp_ln133_29_fu_3277_p2 | icmp_ln133_28_fu_3271_p2);

    assign or_ln133_15_fu_3301_p2 = (icmp_ln133_31_fu_3295_p2 | icmp_ln133_30_fu_3289_p2);

    assign or_ln133_1_fu_1373_p2 = (icmp_ln133_3_fu_1367_p2 | icmp_ln133_2_fu_1361_p2);

    assign or_ln133_2_fu_1564_p2 = (icmp_ln133_5_fu_1558_p2 | icmp_ln133_4_fu_1552_p2);

    assign or_ln133_3_fu_1582_p2 = (icmp_ln133_7_fu_1576_p2 | icmp_ln133_6_fu_1570_p2);

    assign or_ln133_4_fu_1851_p2 = (icmp_ln133_9_fu_1845_p2 | icmp_ln133_8_fu_1839_p2);

    assign or_ln133_5_fu_1869_p2 = (icmp_ln133_11_fu_1863_p2 | icmp_ln133_10_fu_1857_p2);

    assign or_ln133_6_fu_2138_p2 = (icmp_ln133_13_fu_2132_p2 | icmp_ln133_12_fu_2126_p2);

    assign or_ln133_7_fu_2156_p2 = (icmp_ln133_15_fu_2150_p2 | icmp_ln133_14_fu_2144_p2);

    assign or_ln133_8_fu_2422_p2 = (icmp_ln133_17_fu_2416_p2 | icmp_ln133_16_fu_2410_p2);

    assign or_ln133_9_fu_2440_p2 = (icmp_ln133_19_fu_2434_p2 | icmp_ln133_18_fu_2428_p2);

    assign or_ln133_fu_1355_p2 = (icmp_ln133_fu_1343_p2 | icmp_ln133_1_fu_1349_p2);

    assign or_ln134_1_fu_1923_p2 = (icmp_ln134_3_fu_1917_p2 | icmp_ln134_2_fu_1911_p2);

    assign or_ln134_2_fu_2210_p2 = (icmp_ln134_5_fu_2204_p2 | icmp_ln134_4_fu_2198_p2);

    assign or_ln134_3_fu_2494_p2 = (icmp_ln134_7_fu_2488_p2 | icmp_ln134_6_fu_2482_p2);

    assign or_ln134_4_fu_2781_p2 = (icmp_ln134_9_fu_2775_p2 | icmp_ln134_8_fu_2769_p2);

    assign or_ln134_5_fu_3068_p2 = (icmp_ln134_11_fu_3062_p2 | icmp_ln134_10_fu_3056_p2);

    assign or_ln134_6_fu_3355_p2 = (icmp_ln134_13_fu_3349_p2 | icmp_ln134_12_fu_3343_p2);

    assign or_ln134_fu_1636_p2 = (icmp_ln134_fu_1624_p2 | icmp_ln134_1_fu_1630_p2);

    assign or_ln135_10_fu_2853_p2 = (icmp_ln135_21_fu_2847_p2 | icmp_ln135_20_fu_2841_p2);

    assign or_ln135_11_fu_2871_p2 = (icmp_ln135_23_fu_2865_p2 | icmp_ln135_22_fu_2859_p2);

    assign or_ln135_12_fu_3140_p2 = (icmp_ln135_25_fu_3134_p2 | icmp_ln135_24_fu_3128_p2);

    assign or_ln135_13_fu_3158_p2 = (icmp_ln135_27_fu_3152_p2 | icmp_ln135_26_fu_3146_p2);

    assign or_ln135_14_fu_3426_p2 = (icmp_ln135_29_fu_3420_p2 | icmp_ln135_28_fu_3414_p2);

    assign or_ln135_15_fu_3444_p2 = (icmp_ln135_31_fu_3438_p2 | icmp_ln135_30_fu_3432_p2);

    assign or_ln135_1_fu_1479_p2 = (icmp_ln135_3_fu_1473_p2 | icmp_ln135_2_fu_1467_p2);

    assign or_ln135_2_fu_1708_p2 = (icmp_ln135_5_fu_1702_p2 | icmp_ln135_4_fu_1696_p2);

    assign or_ln135_3_fu_1726_p2 = (icmp_ln135_7_fu_1720_p2 | icmp_ln135_6_fu_1714_p2);

    assign or_ln135_4_fu_1995_p2 = (icmp_ln135_9_fu_1989_p2 | icmp_ln135_8_fu_1983_p2);

    assign or_ln135_5_fu_2013_p2 = (icmp_ln135_11_fu_2007_p2 | icmp_ln135_10_fu_2001_p2);

    assign or_ln135_6_fu_2281_p2 = (icmp_ln135_13_fu_2275_p2 | icmp_ln135_12_fu_2269_p2);

    assign or_ln135_7_fu_2299_p2 = (icmp_ln135_15_fu_2293_p2 | icmp_ln135_14_fu_2287_p2);

    assign or_ln135_8_fu_2566_p2 = (icmp_ln135_17_fu_2560_p2 | icmp_ln135_16_fu_2554_p2);

    assign or_ln135_9_fu_2584_p2 = (icmp_ln135_19_fu_2578_p2 | icmp_ln135_18_fu_2572_p2);

    assign or_ln135_fu_1461_p2 = (icmp_ln135_fu_1449_p2 | icmp_ln135_1_fu_1455_p2);

    assign or_ln136_1_fu_2067_p2 = (icmp_ln136_3_fu_2061_p2 | icmp_ln136_2_fu_2055_p2);

    assign or_ln136_2_fu_2352_p2 = (icmp_ln136_5_fu_2346_p2 | icmp_ln136_4_fu_2340_p2);

    assign or_ln136_3_fu_2638_p2 = (icmp_ln136_7_fu_2632_p2 | icmp_ln136_6_fu_2626_p2);

    assign or_ln136_4_fu_2925_p2 = (icmp_ln136_9_fu_2919_p2 | icmp_ln136_8_fu_2913_p2);

    assign or_ln136_5_fu_3212_p2 = (icmp_ln136_11_fu_3206_p2 | icmp_ln136_10_fu_3200_p2);

    assign or_ln136_6_fu_3497_p2 = (icmp_ln136_13_fu_3491_p2 | icmp_ln136_12_fu_3485_p2);

    assign or_ln136_fu_1780_p2 = (icmp_ln136_fu_1768_p2 | icmp_ln136_1_fu_1774_p2);

    assign or_ln139_1_fu_3585_p2 = (icmp_ln139_3_fu_3579_p2 | icmp_ln139_2_fu_3573_p2);

    assign or_ln139_2_fu_3626_p2 = (icmp_ln139_5_fu_3620_p2 | icmp_ln139_4_fu_3614_p2);

    assign or_ln139_fu_3567_p2 = (icmp_ln139_fu_3555_p2 | icmp_ln139_1_fu_3561_p2);

    assign or_ln140_1_fu_3672_p2 = (icmp_ln140_fu_3660_p2 | icmp_ln140_1_fu_3666_p2);

    assign or_ln140_2_fu_3727_p2 = (and_ln142_fu_3722_p2 | and_ln140_reg_5052);

    assign or_ln140_fu_3705_p2 = (and_ln141_fu_3700_p2 | and_ln140_4_fu_3695_p2);

    assign p2_0_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_0_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_0_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_1_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_1_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_1_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_2_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_2_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_2_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_3_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_3_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_3_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_4_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_4_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_4_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_5_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_5_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_5_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_6_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_6_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_6_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_7_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_7_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_7_2_address0 = p2_offset_cast_fu_934_p1;

    assign p2_8_0_address0 = p2_offset_cast_fu_934_p1;

    assign p2_8_1_address0 = p2_offset_cast_fu_934_p1;

    assign p2_8_2_address0 = p2_offset_cast_reg_3746;

    assign p2_offset_cast_fu_934_p1 = p2_offset;

    assign sext_ln120_fu_1001_p1 = $signed(sub_ln120_fu_995_p2);

    assign shl_ln120_fu_1031_p2 = add_ln120_2_reg_3786 << 6'd2;

    assign sub_ln120_1_fu_1036_p2 = (shl_ln120_fu_1031_p2 - add_ln120_2_reg_3786);

    assign sub_ln120_fu_995_p2 = (zext_ln120_5_fu_991_p1 - zext_ln120_fu_964_p1);

    assign tmp_11_fu_1610_p4 = {{bitcast_ln134_fu_1607_p1[62:52]}};

    assign tmp_13_fu_1665_p4 = {{bitcast_ln135_2_fu_1661_p1[62:52]}};

    assign tmp_14_fu_1682_p4 = {{bitcast_ln135_3_fu_1679_p1[62:52]}};

    assign tmp_16_fu_1754_p4 = {{bitcast_ln136_fu_1751_p1[62:52]}};

    assign tmp_18_fu_1808_p4 = {{bitcast_ln133_4_fu_1804_p1[62:52]}};

    assign tmp_19_fu_1825_p4 = {{bitcast_ln133_5_fu_1822_p1[62:52]}};

    assign tmp_1_fu_1311_p4 = {{bitcast_ln133_fu_1307_p1[62:52]}};

    assign tmp_21_fu_1897_p4 = {{bitcast_ln134_1_fu_1894_p1[62:52]}};

    assign tmp_23_fu_1952_p4 = {{bitcast_ln135_4_fu_1948_p1[62:52]}};

    assign tmp_24_fu_1969_p4 = {{bitcast_ln135_5_fu_1966_p1[62:52]}};

    assign tmp_26_fu_2041_p4 = {{bitcast_ln136_1_fu_2038_p1[62:52]}};

    assign tmp_28_fu_2095_p4 = {{bitcast_ln133_6_fu_2091_p1[62:52]}};

    assign tmp_29_fu_2112_p4 = {{bitcast_ln133_7_fu_2109_p1[62:52]}};

    assign tmp_2_fu_1329_p4 = {{bitcast_ln133_1_fu_1325_p1[62:52]}};

    assign tmp_31_fu_2184_p4 = {{bitcast_ln134_2_fu_2181_p1[62:52]}};

    assign tmp_33_fu_2238_p4 = {{bitcast_ln135_6_fu_2235_p1[62:52]}};

    assign tmp_34_fu_2255_p4 = {{bitcast_ln135_7_fu_2252_p1[62:52]}};

    assign tmp_36_fu_2326_p4 = {{bitcast_ln136_2_fu_2323_p1[62:52]}};

    assign tmp_38_fu_2379_p4 = {{bitcast_ln133_8_fu_2375_p1[62:52]}};

    assign tmp_39_fu_2396_p4 = {{bitcast_ln133_9_fu_2393_p1[62:52]}};

    assign tmp_41_fu_2468_p4 = {{bitcast_ln134_3_fu_2465_p1[62:52]}};

    assign tmp_43_fu_2523_p4 = {{bitcast_ln135_8_fu_2519_p1[62:52]}};

    assign tmp_44_fu_2540_p4 = {{bitcast_ln135_9_fu_2537_p1[62:52]}};

    assign tmp_46_fu_2612_p4 = {{bitcast_ln136_3_fu_2609_p1[62:52]}};

    assign tmp_48_fu_2666_p4 = {{bitcast_ln133_10_fu_2662_p1[62:52]}};

    assign tmp_49_fu_2683_p4 = {{bitcast_ln133_11_fu_2680_p1[62:52]}};

    assign tmp_4_fu_1521_p4 = {{bitcast_ln133_2_fu_1517_p1[62:52]}};

    assign tmp_51_fu_2755_p4 = {{bitcast_ln134_4_fu_2752_p1[62:52]}};

    assign tmp_53_fu_2810_p4 = {{bitcast_ln135_10_fu_2806_p1[62:52]}};

    assign tmp_54_fu_2827_p4 = {{bitcast_ln135_11_fu_2824_p1[62:52]}};

    assign tmp_56_fu_2899_p4 = {{bitcast_ln136_4_fu_2896_p1[62:52]}};

    assign tmp_58_fu_2953_p4 = {{bitcast_ln133_12_fu_2949_p1[62:52]}};

    assign tmp_59_fu_2970_p4 = {{bitcast_ln133_13_fu_2967_p1[62:52]}};

    assign tmp_5_fu_1538_p4 = {{bitcast_ln133_3_fu_1535_p1[62:52]}};

    assign tmp_61_fu_3042_p4 = {{bitcast_ln134_5_fu_3039_p1[62:52]}};

    assign tmp_63_fu_3097_p4 = {{bitcast_ln135_12_fu_3093_p1[62:52]}};

    assign tmp_64_fu_3114_p4 = {{bitcast_ln135_13_fu_3111_p1[62:52]}};

    assign tmp_66_fu_3186_p4 = {{bitcast_ln136_5_fu_3183_p1[62:52]}};

    assign tmp_68_fu_3240_p4 = {{bitcast_ln133_14_fu_3236_p1[62:52]}};

    assign tmp_69_fu_3257_p4 = {{bitcast_ln133_15_fu_3254_p1[62:52]}};

    assign tmp_71_fu_3329_p4 = {{bitcast_ln134_6_fu_3326_p1[62:52]}};

    assign tmp_73_fu_3383_p4 = {{bitcast_ln135_14_fu_3380_p1[62:52]}};

    assign tmp_74_fu_3400_p4 = {{bitcast_ln135_15_fu_3397_p1[62:52]}};

    assign tmp_76_fu_3471_p4 = {{bitcast_ln136_6_fu_3468_p1[62:52]}};

    assign tmp_78_fu_3524_p4 = {{bitcast_ln139_fu_3521_p1[62:52]}};

    assign tmp_79_fu_3541_p4 = {{bitcast_ln139_1_fu_3538_p1[62:52]}};

    assign tmp_7_fu_1417_p4 = {{bitcast_ln135_fu_1413_p1[62:52]}};

    assign tmp_81_fu_3600_p4 = {{bitcast_ln139_2_fu_3597_p1[62:52]}};

    assign tmp_83_fu_3646_p4 = {{bitcast_ln140_fu_3643_p1[62:52]}};

    assign tmp_8_fu_1435_p4 = {{bitcast_ln135_1_fu_1431_p1[62:52]}};

    assign tmp_fu_983_p3 = {{p1_offset}, {2'd0}};

    assign trunc_ln133_10_fu_2676_p1 = bitcast_ln133_10_fu_2662_p1[51:0];

    assign trunc_ln133_11_fu_2693_p1 = bitcast_ln133_11_fu_2680_p1[51:0];

    assign trunc_ln133_12_fu_2963_p1 = bitcast_ln133_12_fu_2949_p1[51:0];

    assign trunc_ln133_13_fu_2980_p1 = bitcast_ln133_13_fu_2967_p1[51:0];

    assign trunc_ln133_14_fu_3250_p1 = bitcast_ln133_14_fu_3236_p1[51:0];

    assign trunc_ln133_15_fu_3267_p1 = bitcast_ln133_15_fu_3254_p1[51:0];

    assign trunc_ln133_1_fu_1339_p1 = bitcast_ln133_1_fu_1325_p1[51:0];

    assign trunc_ln133_2_fu_1531_p1 = bitcast_ln133_2_fu_1517_p1[51:0];

    assign trunc_ln133_3_fu_1548_p1 = bitcast_ln133_3_fu_1535_p1[51:0];

    assign trunc_ln133_4_fu_1818_p1 = bitcast_ln133_4_fu_1804_p1[51:0];

    assign trunc_ln133_5_fu_1835_p1 = bitcast_ln133_5_fu_1822_p1[51:0];

    assign trunc_ln133_6_fu_2105_p1 = bitcast_ln133_6_fu_2091_p1[51:0];

    assign trunc_ln133_7_fu_2122_p1 = bitcast_ln133_7_fu_2109_p1[51:0];

    assign trunc_ln133_8_fu_2389_p1 = bitcast_ln133_8_fu_2375_p1[51:0];

    assign trunc_ln133_9_fu_2406_p1 = bitcast_ln133_9_fu_2393_p1[51:0];

    assign trunc_ln133_fu_1321_p1 = bitcast_ln133_fu_1307_p1[51:0];

    assign trunc_ln134_1_fu_1907_p1 = bitcast_ln134_1_fu_1894_p1[51:0];

    assign trunc_ln134_2_fu_2194_p1 = bitcast_ln134_2_fu_2181_p1[51:0];

    assign trunc_ln134_3_fu_2478_p1 = bitcast_ln134_3_fu_2465_p1[51:0];

    assign trunc_ln134_4_fu_2765_p1 = bitcast_ln134_4_fu_2752_p1[51:0];

    assign trunc_ln134_5_fu_3052_p1 = bitcast_ln134_5_fu_3039_p1[51:0];

    assign trunc_ln134_6_fu_3339_p1 = bitcast_ln134_6_fu_3326_p1[51:0];

    assign trunc_ln134_fu_1620_p1 = bitcast_ln134_fu_1607_p1[51:0];

    assign trunc_ln135_10_fu_2820_p1 = bitcast_ln135_10_fu_2806_p1[51:0];

    assign trunc_ln135_11_fu_2837_p1 = bitcast_ln135_11_fu_2824_p1[51:0];

    assign trunc_ln135_12_fu_3107_p1 = bitcast_ln135_12_fu_3093_p1[51:0];

    assign trunc_ln135_13_fu_3124_p1 = bitcast_ln135_13_fu_3111_p1[51:0];

    assign trunc_ln135_14_fu_3393_p1 = bitcast_ln135_14_fu_3380_p1[51:0];

    assign trunc_ln135_15_fu_3410_p1 = bitcast_ln135_15_fu_3397_p1[51:0];

    assign trunc_ln135_1_fu_1445_p1 = bitcast_ln135_1_fu_1431_p1[51:0];

    assign trunc_ln135_2_fu_1675_p1 = bitcast_ln135_2_fu_1661_p1[51:0];

    assign trunc_ln135_3_fu_1692_p1 = bitcast_ln135_3_fu_1679_p1[51:0];

    assign trunc_ln135_4_fu_1962_p1 = bitcast_ln135_4_fu_1948_p1[51:0];

    assign trunc_ln135_5_fu_1979_p1 = bitcast_ln135_5_fu_1966_p1[51:0];

    assign trunc_ln135_6_fu_2248_p1 = bitcast_ln135_6_fu_2235_p1[51:0];

    assign trunc_ln135_7_fu_2265_p1 = bitcast_ln135_7_fu_2252_p1[51:0];

    assign trunc_ln135_8_fu_2533_p1 = bitcast_ln135_8_fu_2519_p1[51:0];

    assign trunc_ln135_9_fu_2550_p1 = bitcast_ln135_9_fu_2537_p1[51:0];

    assign trunc_ln135_fu_1427_p1 = bitcast_ln135_fu_1413_p1[51:0];

    assign trunc_ln136_1_fu_2051_p1 = bitcast_ln136_1_fu_2038_p1[51:0];

    assign trunc_ln136_2_fu_2336_p1 = bitcast_ln136_2_fu_2323_p1[51:0];

    assign trunc_ln136_3_fu_2622_p1 = bitcast_ln136_3_fu_2609_p1[51:0];

    assign trunc_ln136_4_fu_2909_p1 = bitcast_ln136_4_fu_2896_p1[51:0];

    assign trunc_ln136_5_fu_3196_p1 = bitcast_ln136_5_fu_3183_p1[51:0];

    assign trunc_ln136_6_fu_3481_p1 = bitcast_ln136_6_fu_3468_p1[51:0];

    assign trunc_ln136_fu_1764_p1 = bitcast_ln136_fu_1751_p1[51:0];

    assign trunc_ln139_1_fu_3551_p1 = bitcast_ln139_1_fu_3538_p1[51:0];

    assign trunc_ln139_2_fu_3610_p1 = bitcast_ln139_2_fu_3597_p1[51:0];

    assign trunc_ln139_fu_3534_p1 = bitcast_ln139_fu_3521_p1[51:0];

    assign trunc_ln140_fu_3656_p1 = bitcast_ln140_fu_3643_p1[51:0];

    assign zext_ln120_2_fu_978_p1 = mul_ln120_fu_972_p2;

    assign zext_ln120_3_fu_1092_p1 = add_ln120_fu_1087_p2;

    assign zext_ln120_4_fu_1172_p1 = add_ln120_1_fu_1167_p2;

    assign zext_ln120_5_fu_991_p1 = tmp_fu_983_p3;

    assign zext_ln120_6_fu_1041_p1 = sub_ln120_1_fu_1036_p2;

    assign zext_ln120_7_fu_1052_p1 = add_ln120_3_fu_1046_p2;

    assign zext_ln120_8_fu_1082_p1 = add_ln120_4_fu_1077_p2;

    assign zext_ln120_fu_964_p1 = p1_offset;

    assign zext_ln129_10_fu_1152_p1 = add_ln129_10_fu_1147_p2;

    assign zext_ln129_11_fu_1252_p1 = add_ln129_11_fu_1247_p2;

    assign zext_ln129_12_fu_1122_p1 = add_ln129_12_fu_1117_p2;

    assign zext_ln129_13_fu_1192_p1 = add_ln129_13_fu_1187_p2;

    assign zext_ln129_14_fu_1272_p1 = add_ln129_14_fu_1267_p2;

    assign zext_ln129_15_fu_1142_p1 = add_ln129_15_fu_1137_p2;

    assign zext_ln129_16_fu_1222_p1 = add_ln129_16_fu_1217_p2;

    assign zext_ln129_17_fu_1282_p1 = add_ln129_17_fu_1277_p2;

    assign zext_ln129_18_fu_1162_p1 = add_ln129_18_fu_1157_p2;

    assign zext_ln129_19_fu_1242_p1 = add_ln129_19_fu_1237_p2;

    assign zext_ln129_1_fu_1102_p1 = add_ln129_1_fu_1097_p2;

    assign zext_ln129_20_fu_1292_p1 = add_ln129_20_fu_1287_p2;

    assign zext_ln129_21_fu_1202_p1 = add_ln129_21_fu_1197_p2;

    assign zext_ln129_22_fu_1262_p1 = add_ln129_22_fu_1257_p2;

    assign zext_ln129_23_fu_1302_p1 = add_ln129_23_fu_1297_p2;

    assign zext_ln129_2_fu_1182_p1 = add_ln129_2_fu_1177_p2;

    assign zext_ln129_3_fu_1026_p1 = add_ln129_3_fu_1021_p2;

    assign zext_ln129_4_fu_1112_p1 = add_ln129_4_fu_1107_p2;

    assign zext_ln129_5_fu_1212_p1 = add_ln129_5_fu_1207_p2;

    assign zext_ln129_6_fu_1062_p1 = add_ln129_6_fu_1057_p2;

    assign zext_ln129_7_fu_1132_p1 = add_ln129_7_fu_1127_p2;

    assign zext_ln129_8_fu_1232_p1 = add_ln129_8_fu_1227_p2;

    assign zext_ln129_9_fu_1072_p1 = add_ln129_9_fu_1067_p2;

    assign zext_ln129_fu_1016_p1 = add_ln129_fu_1011_p2;

    always @(posedge ap_clk) begin
        p2_offset_cast_reg_3746[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_pointsOverlap_double_2
