/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_pointsOverlap_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    p_read,
    p_read1,
    p_read2,
    ap_return
);

    parameter ap_ST_fsm_pp0_stage0 = 14'd1;
    parameter ap_ST_fsm_pp0_stage1 = 14'd2;
    parameter ap_ST_fsm_pp0_stage2 = 14'd4;
    parameter ap_ST_fsm_pp0_stage3 = 14'd8;
    parameter ap_ST_fsm_pp0_stage4 = 14'd16;
    parameter ap_ST_fsm_pp0_stage5 = 14'd32;
    parameter ap_ST_fsm_pp0_stage6 = 14'd64;
    parameter ap_ST_fsm_pp0_stage7 = 14'd128;
    parameter ap_ST_fsm_pp0_stage8 = 14'd256;
    parameter ap_ST_fsm_pp0_stage9 = 14'd512;
    parameter ap_ST_fsm_pp0_stage10 = 14'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 14'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 14'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 14'd8192;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    input [63:0] p_read;
    input [63:0] p_read1;
    input [63:0] p_read2;
    output [0:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[6:0] p1_address0;
    reg p1_ce0;
    reg[6:0] p1_address1;
    reg p1_ce1;
    reg p2_0_0_ce0;
    reg p2_0_1_ce0;
    reg p2_0_2_ce0;
    reg p2_1_0_ce0;
    reg p2_1_1_ce0;
    reg p2_1_2_ce0;
    reg p2_2_0_ce0;
    reg p2_2_1_ce0;
    reg p2_2_2_ce0;
    reg p2_3_0_ce0;
    reg p2_3_1_ce0;
    reg p2_3_2_ce0;
    reg p2_4_0_ce0;
    reg p2_4_1_ce0;
    reg p2_4_2_ce0;
    reg p2_5_0_ce0;
    reg p2_5_1_ce0;
    reg p2_5_2_ce0;
    reg p2_6_0_ce0;
    reg p2_6_1_ce0;
    reg p2_6_2_ce0;
    reg p2_7_0_ce0;
    reg p2_7_1_ce0;
    reg p2_7_2_ce0;
    reg p2_8_0_ce0;
    reg p2_8_1_ce0;
    reg p2_8_2_ce0;

    (* fsm_encoding = "none" *) reg   [13:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_subdone;
    reg   [63:0] reg_802;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    reg   [63:0] reg_807;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    reg   [63:0] reg_814;
    reg   [63:0] reg_821;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    reg   [63:0] reg_827;
    reg   [63:0] reg_833;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    reg   [63:0] reg_838;
    reg   [63:0] reg_844;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    reg   [63:0] reg_849;
    reg   [63:0] reg_855;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    wire    ap_block_pp0_stage13_11001;
    reg   [63:0] reg_860;
    reg   [63:0] reg_866;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] reg_872;
    wire   [63:0] grp_fu_751_p2;
    reg   [63:0] reg_878;
    wire   [63:0] grp_fu_756_p2;
    reg   [63:0] reg_884;
    wire   [63:0] grp_fu_761_p2;
    reg   [63:0] reg_891;
    reg   [63:0] reg_898;
    reg   [63:0] reg_904;
    reg   [63:0] reg_911;
    reg   [63:0] reg_918;
    reg   [63:0] reg_924;
    reg   [63:0] reg_930;
    reg   [63:0] reg_938;
    reg   [63:0] reg_944;
    wire   [6:0] mul_ln120_fu_984_p2;
    reg   [6:0] mul_ln120_reg_3688;
    reg   [63:0] p2_0_0_load_reg_3868;
    reg   [63:0] p2_0_1_load_reg_3873;
    reg   [63:0] p2_0_2_load_reg_3878;
    reg   [63:0] p2_1_0_load_reg_3883;
    reg   [63:0] p2_1_1_load_reg_3888;
    reg   [63:0] p2_1_2_load_reg_3893;
    reg   [63:0] p2_2_0_load_reg_3898;
    reg   [63:0] p2_2_1_load_reg_3903;
    reg   [63:0] p2_2_2_load_reg_3908;
    reg   [63:0] p2_3_0_load_reg_3913;
    reg   [63:0] p2_3_1_load_reg_3918;
    reg   [63:0] p2_3_2_load_reg_3923;
    reg   [63:0] p2_4_0_load_reg_3928;
    reg   [63:0] p2_4_1_load_reg_3933;
    reg   [63:0] p2_4_2_load_reg_3938;
    reg   [63:0] p2_5_0_load_reg_3943;
    reg   [63:0] p2_5_1_load_reg_3948;
    reg   [63:0] p2_5_2_load_reg_3953;
    reg   [63:0] p2_6_0_load_reg_3958;
    reg   [63:0] p2_6_1_load_reg_3963;
    reg   [63:0] p2_6_2_load_reg_3968;
    reg   [63:0] p2_7_0_load_reg_3973;
    reg   [63:0] p2_7_1_load_reg_3978;
    reg   [63:0] p2_7_2_load_reg_3983;
    reg   [63:0] p2_8_0_load_reg_3988;
    reg   [63:0] p2_8_1_load_reg_3993;
    reg   [63:0] p2_8_2_load_reg_3998;
    reg   [63:0] p_read83_reg_4003;
    reg   [63:0] p_read_65_reg_4031;
    reg   [63:0] p_read_64_reg_4079;
    wire   [63:0] grp_fu_766_p2;
    reg   [63:0] mul_reg_4097;
    wire   [63:0] grp_fu_771_p2;
    reg   [63:0] mul6_reg_4102;
    wire   [63:0] grp_fu_776_p2;
    reg   [63:0] mul2_reg_4107;
    reg   [63:0] p1_load_5_reg_4112;
    wire   [63:0] grp_fu_781_p2;
    reg   [63:0] mul25_1_reg_4117;
    reg   [63:0] mul1_reg_4132;
    reg   [63:0] mul20_1_reg_4137;
    reg   [63:0] mul25_2_reg_4142;
    reg   [63:0] mul25_3_reg_4147;
    reg   [63:0] mul6_1_reg_4162;
    reg   [63:0] mul25_s_reg_4167;
    reg   [63:0] mul20_2_reg_4172;
    reg   [63:0] mul20_3_reg_4177;
    reg   [63:0] mul_1_reg_4192;
    reg   [63:0] mul20_s_reg_4197;
    reg   [63:0] mul25_1_1_reg_4202;
    reg   [63:0] mul25_4_reg_4207;
    reg   [63:0] mul20_1_1_reg_4222;
    reg   [63:0] mul25_2_1_reg_4227;
    reg   [63:0] mul20_4_reg_4232;
    reg   [63:0] mul25_5_reg_4237;
    reg   [63:0] mul20_2_1_reg_4252;
    reg   [63:0] mul25_3_1_reg_4257;
    reg   [63:0] mul20_5_reg_4262;
    reg   [63:0] mul25_6_reg_4267;
    reg   [63:0] mul6_2_reg_4272;
    reg   [63:0] mul25_8_reg_4277;
    reg   [63:0] mul20_3_1_reg_4282;
    reg   [63:0] mul20_6_reg_4287;
    wire   [63:0] grp_fu_746_p2;
    reg   [63:0] max1_33_reg_4292;
    reg   [63:0] mul_2_reg_4297;
    reg   [63:0] mul20_8_reg_4302;
    reg   [63:0] n2_3_reg_4307;
    reg   [63:0] mul25_4_1_reg_4312;
    reg   [63:0] mul25_7_reg_4317;
    reg   [63:0] n1_reg_4322;
    reg   [63:0] n1_3_reg_4327;
    reg   [63:0] mul25_1_2_reg_4332;
    reg   [63:0] n2_6_reg_4337;
    reg   [63:0] mul20_4_1_reg_4342;
    reg   [63:0] mul25_5_1_reg_4347;
    reg   [63:0] mul20_7_reg_4352;
    reg   [63:0] mul20_1_2_reg_4357;
    reg   [63:0] n1_6_reg_4362;
    reg   [63:0] mul25_2_2_reg_4367;
    reg   [63:0] n1_9_reg_4372;
    reg   [63:0] mul20_5_1_reg_4377;
    reg   [63:0] mul25_6_1_reg_4382;
    reg   [63:0] mul20_2_2_reg_4387;
    reg   [63:0] mul25_3_2_reg_4392;
    reg   [63:0] n2_40_reg_4397;
    reg   [63:0] mul20_6_1_reg_4402;
    reg   [63:0] mul25_7_1_reg_4407;
    reg   [63:0] mul20_3_2_reg_4412;
    reg   [63:0] n1_40_reg_4417;
    reg   [63:0] mul25_4_2_reg_4422;
    reg   [63:0] n2_43_reg_4427;
    reg   [63:0] mul25_5_2_reg_4432;
    reg   [63:0] mul20_7_1_reg_4437;
    reg   [63:0] mul20_4_2_reg_4442;
    reg   [63:0] n1_43_reg_4447;
    reg   [63:0] mul20_5_2_reg_4452;
    reg   [63:0] n2_46_reg_4457;
    reg   [63:0] mul25_6_2_reg_4462;
    reg   [63:0] mul25_7_2_reg_4467;
    reg   [63:0] mul25_7_2_reg_4467_pp0_iter2_reg;
    reg   [63:0] n1_46_reg_4472;
    reg   [63:0] mul20_6_2_reg_4477;
    reg   [63:0] mul20_7_2_reg_4482;
    reg   [63:0] mul20_7_2_reg_4482_pp0_iter2_reg;
    reg   [63:0] max1_1_reg_4487;
    reg   [63:0] n1_1_reg_4492;
    reg   [63:0] n1_4_reg_4497;
    reg   [63:0] n2_38_reg_4502;
    reg   [63:0] n1_7_reg_4507;
    reg   [63:0] n1_38_reg_4512;
    reg   [63:0] n1_49_reg_4517;
    reg   [63:0] n2_49_reg_4522;
    reg   [63:0] n2_41_reg_4527;
    reg   [63:0] n1_41_reg_4532;
    reg   [63:0] n2_44_reg_4537;
    reg   [63:0] n1_44_reg_4542;
    reg   [63:0] n2_47_reg_4547;
    reg   [63:0] n1_47_reg_4552;
    wire   [0:0] and_ln133_fu_1327_p2;
    reg   [0:0] and_ln133_reg_4557;
    wire   [0:0] grp_fu_790_p2;
    reg   [0:0] tmp_176_reg_4563;
    wire   [63:0] max2_fu_1417_p3;
    reg   [63:0] max2_reg_4568;
    wire   [63:0] min2_20_fu_1431_p3;
    reg   [63:0] min2_20_reg_4575;
    wire   [63:0] max1_fu_1443_p3;
    reg   [63:0] max1_reg_4582;
    wire   [63:0] min1_20_fu_1457_p3;
    reg   [63:0] min1_20_reg_4589;
    reg   [63:0] n1_39_reg_4596;
    reg   [63:0] n2_50_reg_4604;
    wire   [0:0] or_ln133_32_fu_1512_p2;
    reg   [0:0] or_ln133_32_reg_4609;
    wire   [63:0] max1_26_fu_1548_p3;
    reg   [63:0] max1_26_reg_4614;
    wire   [63:0] max2_26_fu_1638_p3;
    reg   [63:0] max2_26_reg_4621;
    wire   [63:0] min2_21_fu_1692_p3;
    reg   [63:0] min2_21_reg_4628;
    wire   [63:0] min1_21_fu_1745_p3;
    reg   [63:0] min1_21_reg_4635;
    wire   [0:0] or_ln133_34_fu_1799_p2;
    reg   [0:0] or_ln133_34_reg_4642;
    wire   [63:0] max1_27_fu_1835_p3;
    reg   [63:0] max1_27_reg_4647;
    wire   [63:0] max2_27_fu_1925_p3;
    reg   [63:0] max2_27_reg_4654;
    wire   [63:0] min2_22_fu_1979_p3;
    reg   [63:0] min2_22_reg_4661;
    wire   [63:0] min1_22_fu_2032_p3;
    reg   [63:0] min1_22_reg_4668;
    wire   [0:0] or_ln133_36_fu_2085_p2;
    reg   [0:0] or_ln133_36_reg_4675;
    wire   [63:0] max1_28_fu_2121_p3;
    reg   [63:0] max1_28_reg_4680;
    wire   [63:0] max2_28_fu_2210_p3;
    reg   [63:0] max2_28_reg_4687;
    wire   [63:0] min2_23_fu_2264_p3;
    reg   [63:0] min2_23_reg_4694;
    wire   [63:0] min1_23_fu_2317_p3;
    reg   [63:0] min1_23_reg_4701;
    reg   [63:0] n1_48_reg_4708;
    wire   [0:0] or_ln133_38_fu_2370_p2;
    reg   [0:0] or_ln133_38_reg_4716;
    wire   [63:0] max1_29_fu_2406_p3;
    reg   [63:0] max1_29_reg_4721;
    wire   [63:0] max2_29_fu_2496_p3;
    reg   [63:0] max2_29_reg_4728;
    wire   [63:0] min2_24_fu_2550_p3;
    reg   [63:0] min2_24_reg_4735;
    reg   [63:0] n1_51_reg_4742;
    reg   [63:0] n2_51_reg_4751;
    wire   [63:0] min1_24_fu_2603_p3;
    reg   [63:0] min1_24_reg_4760;
    wire   [0:0] or_ln133_40_fu_2657_p2;
    reg   [0:0] or_ln133_40_reg_4767;
    wire   [63:0] max1_30_fu_2693_p3;
    reg   [63:0] max1_30_reg_4772;
    wire   [63:0] max2_30_fu_2783_p3;
    reg   [63:0] max2_30_reg_4779;
    wire   [63:0] min2_25_fu_2837_p3;
    reg   [63:0] min2_25_reg_4786;
    wire   [63:0] min1_25_fu_2890_p3;
    reg   [63:0] min1_25_reg_4793;
    wire   [0:0] or_ln133_42_fu_2943_p2;
    reg   [0:0] or_ln133_42_reg_4800;
    wire   [63:0] max1_31_fu_2979_p3;
    reg   [63:0] max1_31_reg_4805;
    wire   [63:0] max2_31_fu_3068_p3;
    reg   [63:0] max2_31_reg_4812;
    wire   [63:0] min2_26_fu_3122_p3;
    reg   [63:0] min2_26_reg_4819;
    wire   [63:0] min1_26_fu_3175_p3;
    reg   [63:0] min1_26_reg_4826;
    wire   [63:0] max2_32_fu_3263_p3;
    reg   [63:0] max2_32_reg_4833;
    wire   [63:0] min2_27_fu_3316_p3;
    reg   [63:0] min2_27_reg_4841;
    wire   [63:0] max1_32_fu_3404_p3;
    reg   [63:0] max1_32_reg_4848;
    wire   [63:0] min1_27_fu_3457_p3;
    reg   [63:0] min1_27_reg_4855;
    wire   [0:0] grp_fu_794_p2;
    reg   [0:0] tmp_256_reg_4863;
    wire   [0:0] grp_fu_798_p2;
    reg   [0:0] tmp_258_reg_4868;
    reg   [0:0] tmp_259_reg_4873;
    reg   [0:0] tmp_260_reg_4878;
    wire   [0:0] and_ln139_9_fu_3533_p2;
    reg   [0:0] and_ln139_9_reg_4883;
    wire   [0:0] and_ln139_12_fu_3580_p2;
    reg   [0:0] and_ln139_12_reg_4888;
    wire   [0:0] and_ln140_11_fu_3631_p2;
    reg   [0:0] and_ln140_11_reg_4894;
    wire   [0:0] and_ln140_fu_3653_p2;
    reg   [0:0] and_ln140_reg_4899;
    reg   [0:0] tmp_254_reg_4904;
    wire   [0:0] or_ln140_8_fu_3669_p2;
    reg   [0:0] or_ln140_8_reg_4909;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage2_subdone;
    reg   [63:0] ap_port_reg_p_read;
    reg   [63:0] ap_port_reg_p_read1;
    reg   [63:0] ap_port_reg_p_read2;
    wire   [63:0] zext_ln120_17_fu_990_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] p2_offset_cast_fu_949_p1;
    wire   [63:0] zext_ln129_fu_1000_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln129_49_fu_1010_p1;
    wire   [63:0] zext_ln129_52_fu_1020_p1;
    wire    ap_block_pp0_stage2;
    wire   [63:0] zext_ln129_55_fu_1030_p1;
    wire   [63:0] zext_ln120_18_fu_1040_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln129_47_fu_1050_p1;
    wire   [63:0] zext_ln129_50_fu_1060_p1;
    wire    ap_block_pp0_stage4;
    wire   [63:0] zext_ln129_58_fu_1070_p1;
    wire   [63:0] zext_ln129_53_fu_1080_p1;
    wire    ap_block_pp0_stage5;
    wire   [63:0] zext_ln129_61_fu_1090_p1;
    wire   [63:0] zext_ln129_56_fu_1100_p1;
    wire    ap_block_pp0_stage6;
    wire   [63:0] zext_ln129_64_fu_1110_p1;
    wire   [63:0] zext_ln120_19_fu_1120_p1;
    wire    ap_block_pp0_stage7;
    wire   [63:0] zext_ln129_48_fu_1130_p1;
    wire   [63:0] zext_ln129_59_fu_1140_p1;
    wire    ap_block_pp0_stage8;
    wire   [63:0] zext_ln129_67_fu_1150_p1;
    wire   [63:0] zext_ln129_51_fu_1160_p1;
    wire    ap_block_pp0_stage9;
    wire   [63:0] zext_ln129_62_fu_1170_p1;
    wire   [63:0] zext_ln129_54_fu_1180_p1;
    wire    ap_block_pp0_stage10;
    wire   [63:0] zext_ln129_65_fu_1190_p1;
    wire   [63:0] zext_ln129_57_fu_1200_p1;
    wire    ap_block_pp0_stage11;
    wire   [63:0] zext_ln129_68_fu_1210_p1;
    wire   [63:0] zext_ln129_60_fu_1220_p1;
    wire    ap_block_pp0_stage12;
    wire   [63:0] zext_ln129_63_fu_1230_p1;
    wire   [63:0] zext_ln129_66_fu_1240_p1;
    wire    ap_block_pp0_stage13;
    wire   [63:0] zext_ln129_69_fu_1250_p1;
    reg   [63:0] grp_fu_746_p0;
    reg   [63:0] grp_fu_746_p1;
    reg   [63:0] grp_fu_751_p0;
    reg   [63:0] grp_fu_751_p1;
    reg   [63:0] grp_fu_756_p0;
    reg   [63:0] grp_fu_756_p1;
    reg   [63:0] grp_fu_761_p0;
    reg   [63:0] grp_fu_761_p1;
    reg   [63:0] grp_fu_766_p0;
    reg   [63:0] grp_fu_766_p1;
    reg   [63:0] grp_fu_771_p0;
    reg   [63:0] grp_fu_771_p1;
    reg   [63:0] grp_fu_776_p0;
    reg   [63:0] grp_fu_776_p1;
    reg   [63:0] grp_fu_781_p0;
    reg   [63:0] grp_fu_781_p1;
    reg   [63:0] grp_fu_790_p0;
    reg   [63:0] grp_fu_790_p1;
    reg   [63:0] grp_fu_794_p0;
    reg   [63:0] grp_fu_794_p1;
    reg   [63:0] grp_fu_798_p0;
    reg   [63:0] grp_fu_798_p1;
    wire   [1:0] mul_ln120_fu_984_p0;
    wire   [5:0] mul_ln120_fu_984_p1;
    wire   [6:0] add_ln129_fu_995_p2;
    wire   [6:0] add_ln129_49_fu_1005_p2;
    wire   [6:0] add_ln129_52_fu_1015_p2;
    wire   [6:0] add_ln129_55_fu_1025_p2;
    wire   [6:0] add_ln120_fu_1035_p2;
    wire   [6:0] add_ln129_47_fu_1045_p2;
    wire   [6:0] add_ln129_50_fu_1055_p2;
    wire   [6:0] add_ln129_58_fu_1065_p2;
    wire   [6:0] add_ln129_53_fu_1075_p2;
    wire   [6:0] add_ln129_61_fu_1085_p2;
    wire   [6:0] add_ln129_56_fu_1095_p2;
    wire   [6:0] add_ln129_64_fu_1105_p2;
    wire   [6:0] add_ln120_9_fu_1115_p2;
    wire   [6:0] add_ln129_48_fu_1125_p2;
    wire   [6:0] add_ln129_59_fu_1135_p2;
    wire   [6:0] add_ln129_67_fu_1145_p2;
    wire   [6:0] add_ln129_51_fu_1155_p2;
    wire   [6:0] add_ln129_62_fu_1165_p2;
    wire   [6:0] add_ln129_54_fu_1175_p2;
    wire   [6:0] add_ln129_65_fu_1185_p2;
    wire   [6:0] add_ln129_57_fu_1195_p2;
    wire   [6:0] add_ln129_68_fu_1205_p2;
    wire   [6:0] add_ln129_60_fu_1215_p2;
    wire   [6:0] add_ln129_63_fu_1225_p2;
    wire   [6:0] add_ln129_66_fu_1235_p2;
    wire   [6:0] add_ln129_69_fu_1245_p2;
    wire   [63:0] bitcast_ln133_fu_1255_p1;
    wire   [63:0] bitcast_ln133_31_fu_1273_p1;
    wire   [10:0] tmp_s_fu_1259_p4;
    wire   [51:0] trunc_ln133_fu_1269_p1;
    wire   [0:0] icmp_ln133_63_fu_1297_p2;
    wire   [0:0] icmp_ln133_fu_1291_p2;
    wire   [10:0] tmp_175_fu_1277_p4;
    wire   [51:0] trunc_ln133_31_fu_1287_p1;
    wire   [0:0] icmp_ln133_65_fu_1315_p2;
    wire   [0:0] icmp_ln133_64_fu_1309_p2;
    wire   [0:0] or_ln133_fu_1303_p2;
    wire   [0:0] or_ln133_31_fu_1321_p2;
    wire   [63:0] bitcast_ln135_fu_1333_p1;
    wire   [63:0] bitcast_ln135_31_fu_1351_p1;
    wire   [10:0] tmp_178_fu_1337_p4;
    wire   [51:0] trunc_ln135_fu_1347_p1;
    wire   [0:0] icmp_ln135_63_fu_1375_p2;
    wire   [0:0] icmp_ln135_fu_1369_p2;
    wire   [10:0] tmp_179_fu_1355_p4;
    wire   [51:0] trunc_ln135_31_fu_1365_p1;
    wire   [0:0] icmp_ln135_65_fu_1393_p2;
    wire   [0:0] icmp_ln135_64_fu_1387_p2;
    wire   [0:0] or_ln135_fu_1381_p2;
    wire   [0:0] or_ln135_31_fu_1399_p2;
    wire   [0:0] and_ln135_fu_1405_p2;
    wire   [0:0] and_ln135_31_fu_1411_p2;
    wire   [0:0] and_ln136_fu_1425_p2;
    wire   [0:0] and_ln133_31_fu_1439_p2;
    wire   [0:0] and_ln134_fu_1452_p2;
    wire   [63:0] bitcast_ln133_32_fu_1465_p1;
    wire   [63:0] bitcast_ln133_33_fu_1483_p1;
    wire   [10:0] tmp_182_fu_1469_p4;
    wire   [51:0] trunc_ln133_32_fu_1479_p1;
    wire   [0:0] icmp_ln133_67_fu_1506_p2;
    wire   [0:0] icmp_ln133_66_fu_1500_p2;
    wire   [10:0] tmp_183_fu_1486_p4;
    wire   [51:0] trunc_ln133_33_fu_1496_p1;
    wire   [0:0] icmp_ln133_69_fu_1524_p2;
    wire   [0:0] icmp_ln133_68_fu_1518_p2;
    wire   [0:0] or_ln133_33_fu_1530_p2;
    wire   [0:0] and_ln133_32_fu_1536_p2;
    wire   [0:0] and_ln133_33_fu_1542_p2;
    wire   [63:0] bitcast_ln135_32_fu_1555_p1;
    wire   [63:0] bitcast_ln135_33_fu_1573_p1;
    wire   [10:0] tmp_187_fu_1559_p4;
    wire   [51:0] trunc_ln135_32_fu_1569_p1;
    wire   [0:0] icmp_ln135_67_fu_1596_p2;
    wire   [0:0] icmp_ln135_66_fu_1590_p2;
    wire   [10:0] tmp_188_fu_1576_p4;
    wire   [51:0] trunc_ln135_33_fu_1586_p1;
    wire   [0:0] icmp_ln135_69_fu_1614_p2;
    wire   [0:0] icmp_ln135_68_fu_1608_p2;
    wire   [0:0] or_ln135_32_fu_1602_p2;
    wire   [0:0] or_ln135_33_fu_1620_p2;
    wire   [0:0] and_ln135_32_fu_1626_p2;
    wire   [0:0] and_ln135_33_fu_1632_p2;
    wire   [63:0] bitcast_ln136_fu_1645_p1;
    wire   [10:0] tmp_190_fu_1648_p4;
    wire   [51:0] trunc_ln136_fu_1658_p1;
    wire   [0:0] icmp_ln136_27_fu_1668_p2;
    wire   [0:0] icmp_ln136_fu_1662_p2;
    wire   [0:0] or_ln136_fu_1674_p2;
    wire   [0:0] and_ln136_29_fu_1680_p2;
    wire   [0:0] and_ln136_30_fu_1686_p2;
    wire   [63:0] bitcast_ln134_fu_1699_p1;
    wire   [10:0] tmp_185_fu_1702_p4;
    wire   [51:0] trunc_ln134_fu_1712_p1;
    wire   [0:0] icmp_ln134_27_fu_1722_p2;
    wire   [0:0] icmp_ln134_fu_1716_p2;
    wire   [0:0] or_ln134_fu_1728_p2;
    wire   [0:0] and_ln134_29_fu_1734_p2;
    wire   [0:0] and_ln134_30_fu_1739_p2;
    wire   [63:0] bitcast_ln133_34_fu_1752_p1;
    wire   [63:0] bitcast_ln133_35_fu_1770_p1;
    wire   [10:0] tmp_192_fu_1756_p4;
    wire   [51:0] trunc_ln133_34_fu_1766_p1;
    wire   [0:0] icmp_ln133_71_fu_1793_p2;
    wire   [0:0] icmp_ln133_70_fu_1787_p2;
    wire   [10:0] tmp_193_fu_1773_p4;
    wire   [51:0] trunc_ln133_35_fu_1783_p1;
    wire   [0:0] icmp_ln133_73_fu_1811_p2;
    wire   [0:0] icmp_ln133_72_fu_1805_p2;
    wire   [0:0] or_ln133_35_fu_1817_p2;
    wire   [0:0] and_ln133_34_fu_1823_p2;
    wire   [0:0] and_ln133_35_fu_1829_p2;
    wire   [63:0] bitcast_ln135_34_fu_1842_p1;
    wire   [63:0] bitcast_ln135_35_fu_1860_p1;
    wire   [10:0] tmp_197_fu_1846_p4;
    wire   [51:0] trunc_ln135_34_fu_1856_p1;
    wire   [0:0] icmp_ln135_71_fu_1883_p2;
    wire   [0:0] icmp_ln135_70_fu_1877_p2;
    wire   [10:0] tmp_198_fu_1863_p4;
    wire   [51:0] trunc_ln135_35_fu_1873_p1;
    wire   [0:0] icmp_ln135_73_fu_1901_p2;
    wire   [0:0] icmp_ln135_72_fu_1895_p2;
    wire   [0:0] or_ln135_34_fu_1889_p2;
    wire   [0:0] or_ln135_35_fu_1907_p2;
    wire   [0:0] and_ln135_34_fu_1913_p2;
    wire   [0:0] and_ln135_35_fu_1919_p2;
    wire   [63:0] bitcast_ln136_13_fu_1932_p1;
    wire   [10:0] tmp_200_fu_1935_p4;
    wire   [51:0] trunc_ln136_13_fu_1945_p1;
    wire   [0:0] icmp_ln136_29_fu_1955_p2;
    wire   [0:0] icmp_ln136_28_fu_1949_p2;
    wire   [0:0] or_ln136_13_fu_1961_p2;
    wire   [0:0] and_ln136_31_fu_1967_p2;
    wire   [0:0] and_ln136_32_fu_1973_p2;
    wire   [63:0] bitcast_ln134_13_fu_1986_p1;
    wire   [10:0] tmp_195_fu_1989_p4;
    wire   [51:0] trunc_ln134_13_fu_1999_p1;
    wire   [0:0] icmp_ln134_29_fu_2009_p2;
    wire   [0:0] icmp_ln134_28_fu_2003_p2;
    wire   [0:0] or_ln134_13_fu_2015_p2;
    wire   [0:0] and_ln134_31_fu_2021_p2;
    wire   [0:0] and_ln134_32_fu_2026_p2;
    wire   [63:0] bitcast_ln133_36_fu_2039_p1;
    wire   [63:0] bitcast_ln133_37_fu_2056_p1;
    wire   [10:0] tmp_202_fu_2042_p4;
    wire   [51:0] trunc_ln133_36_fu_2052_p1;
    wire   [0:0] icmp_ln133_75_fu_2079_p2;
    wire   [0:0] icmp_ln133_74_fu_2073_p2;
    wire   [10:0] tmp_203_fu_2059_p4;
    wire   [51:0] trunc_ln133_37_fu_2069_p1;
    wire   [0:0] icmp_ln133_77_fu_2097_p2;
    wire   [0:0] icmp_ln133_76_fu_2091_p2;
    wire   [0:0] or_ln133_37_fu_2103_p2;
    wire   [0:0] and_ln133_36_fu_2109_p2;
    wire   [0:0] and_ln133_37_fu_2115_p2;
    wire   [63:0] bitcast_ln135_36_fu_2127_p1;
    wire   [63:0] bitcast_ln135_37_fu_2145_p1;
    wire   [10:0] tmp_207_fu_2131_p4;
    wire   [51:0] trunc_ln135_36_fu_2141_p1;
    wire   [0:0] icmp_ln135_75_fu_2168_p2;
    wire   [0:0] icmp_ln135_74_fu_2162_p2;
    wire   [10:0] tmp_208_fu_2148_p4;
    wire   [51:0] trunc_ln135_37_fu_2158_p1;
    wire   [0:0] icmp_ln135_77_fu_2186_p2;
    wire   [0:0] icmp_ln135_76_fu_2180_p2;
    wire   [0:0] or_ln135_36_fu_2174_p2;
    wire   [0:0] or_ln135_37_fu_2192_p2;
    wire   [0:0] and_ln135_36_fu_2198_p2;
    wire   [0:0] and_ln135_37_fu_2204_p2;
    wire   [63:0] bitcast_ln136_14_fu_2217_p1;
    wire   [10:0] tmp_210_fu_2220_p4;
    wire   [51:0] trunc_ln136_14_fu_2230_p1;
    wire   [0:0] icmp_ln136_31_fu_2240_p2;
    wire   [0:0] icmp_ln136_30_fu_2234_p2;
    wire   [0:0] or_ln136_14_fu_2246_p2;
    wire   [0:0] and_ln136_33_fu_2252_p2;
    wire   [0:0] and_ln136_34_fu_2258_p2;
    wire   [63:0] bitcast_ln134_14_fu_2271_p1;
    wire   [10:0] tmp_205_fu_2274_p4;
    wire   [51:0] trunc_ln134_14_fu_2284_p1;
    wire   [0:0] icmp_ln134_31_fu_2294_p2;
    wire   [0:0] icmp_ln134_30_fu_2288_p2;
    wire   [0:0] or_ln134_14_fu_2300_p2;
    wire   [0:0] and_ln134_33_fu_2306_p2;
    wire   [0:0] and_ln134_34_fu_2311_p2;
    wire   [63:0] bitcast_ln133_38_fu_2323_p1;
    wire   [63:0] bitcast_ln133_39_fu_2341_p1;
    wire   [10:0] tmp_212_fu_2327_p4;
    wire   [51:0] trunc_ln133_38_fu_2337_p1;
    wire   [0:0] icmp_ln133_79_fu_2364_p2;
    wire   [0:0] icmp_ln133_78_fu_2358_p2;
    wire   [10:0] tmp_213_fu_2344_p4;
    wire   [51:0] trunc_ln133_39_fu_2354_p1;
    wire   [0:0] icmp_ln133_81_fu_2382_p2;
    wire   [0:0] icmp_ln133_80_fu_2376_p2;
    wire   [0:0] or_ln133_39_fu_2388_p2;
    wire   [0:0] and_ln133_38_fu_2394_p2;
    wire   [0:0] and_ln133_39_fu_2400_p2;
    wire   [63:0] bitcast_ln135_38_fu_2413_p1;
    wire   [63:0] bitcast_ln135_39_fu_2431_p1;
    wire   [10:0] tmp_217_fu_2417_p4;
    wire   [51:0] trunc_ln135_38_fu_2427_p1;
    wire   [0:0] icmp_ln135_79_fu_2454_p2;
    wire   [0:0] icmp_ln135_78_fu_2448_p2;
    wire   [10:0] tmp_218_fu_2434_p4;
    wire   [51:0] trunc_ln135_39_fu_2444_p1;
    wire   [0:0] icmp_ln135_81_fu_2472_p2;
    wire   [0:0] icmp_ln135_80_fu_2466_p2;
    wire   [0:0] or_ln135_38_fu_2460_p2;
    wire   [0:0] or_ln135_39_fu_2478_p2;
    wire   [0:0] and_ln135_38_fu_2484_p2;
    wire   [0:0] and_ln135_39_fu_2490_p2;
    wire   [63:0] bitcast_ln136_15_fu_2503_p1;
    wire   [10:0] tmp_220_fu_2506_p4;
    wire   [51:0] trunc_ln136_15_fu_2516_p1;
    wire   [0:0] icmp_ln136_33_fu_2526_p2;
    wire   [0:0] icmp_ln136_32_fu_2520_p2;
    wire   [0:0] or_ln136_15_fu_2532_p2;
    wire   [0:0] and_ln136_35_fu_2538_p2;
    wire   [0:0] and_ln136_36_fu_2544_p2;
    wire   [63:0] bitcast_ln134_15_fu_2557_p1;
    wire   [10:0] tmp_215_fu_2560_p4;
    wire   [51:0] trunc_ln134_15_fu_2570_p1;
    wire   [0:0] icmp_ln134_33_fu_2580_p2;
    wire   [0:0] icmp_ln134_32_fu_2574_p2;
    wire   [0:0] or_ln134_15_fu_2586_p2;
    wire   [0:0] and_ln134_35_fu_2592_p2;
    wire   [0:0] and_ln134_36_fu_2597_p2;
    wire   [63:0] bitcast_ln133_40_fu_2610_p1;
    wire   [63:0] bitcast_ln133_41_fu_2628_p1;
    wire   [10:0] tmp_222_fu_2614_p4;
    wire   [51:0] trunc_ln133_40_fu_2624_p1;
    wire   [0:0] icmp_ln133_83_fu_2651_p2;
    wire   [0:0] icmp_ln133_82_fu_2645_p2;
    wire   [10:0] tmp_223_fu_2631_p4;
    wire   [51:0] trunc_ln133_41_fu_2641_p1;
    wire   [0:0] icmp_ln133_85_fu_2669_p2;
    wire   [0:0] icmp_ln133_84_fu_2663_p2;
    wire   [0:0] or_ln133_41_fu_2675_p2;
    wire   [0:0] and_ln133_40_fu_2681_p2;
    wire   [0:0] and_ln133_41_fu_2687_p2;
    wire   [63:0] bitcast_ln135_40_fu_2700_p1;
    wire   [63:0] bitcast_ln135_41_fu_2718_p1;
    wire   [10:0] tmp_227_fu_2704_p4;
    wire   [51:0] trunc_ln135_40_fu_2714_p1;
    wire   [0:0] icmp_ln135_83_fu_2741_p2;
    wire   [0:0] icmp_ln135_82_fu_2735_p2;
    wire   [10:0] tmp_228_fu_2721_p4;
    wire   [51:0] trunc_ln135_41_fu_2731_p1;
    wire   [0:0] icmp_ln135_85_fu_2759_p2;
    wire   [0:0] icmp_ln135_84_fu_2753_p2;
    wire   [0:0] or_ln135_40_fu_2747_p2;
    wire   [0:0] or_ln135_41_fu_2765_p2;
    wire   [0:0] and_ln135_40_fu_2771_p2;
    wire   [0:0] and_ln135_41_fu_2777_p2;
    wire   [63:0] bitcast_ln136_16_fu_2790_p1;
    wire   [10:0] tmp_230_fu_2793_p4;
    wire   [51:0] trunc_ln136_16_fu_2803_p1;
    wire   [0:0] icmp_ln136_35_fu_2813_p2;
    wire   [0:0] icmp_ln136_34_fu_2807_p2;
    wire   [0:0] or_ln136_16_fu_2819_p2;
    wire   [0:0] and_ln136_37_fu_2825_p2;
    wire   [0:0] and_ln136_38_fu_2831_p2;
    wire   [63:0] bitcast_ln134_16_fu_2844_p1;
    wire   [10:0] tmp_225_fu_2847_p4;
    wire   [51:0] trunc_ln134_16_fu_2857_p1;
    wire   [0:0] icmp_ln134_35_fu_2867_p2;
    wire   [0:0] icmp_ln134_34_fu_2861_p2;
    wire   [0:0] or_ln134_16_fu_2873_p2;
    wire   [0:0] and_ln134_37_fu_2879_p2;
    wire   [0:0] and_ln134_38_fu_2884_p2;
    wire   [63:0] bitcast_ln133_42_fu_2897_p1;
    wire   [63:0] bitcast_ln133_43_fu_2914_p1;
    wire   [10:0] tmp_232_fu_2900_p4;
    wire   [51:0] trunc_ln133_42_fu_2910_p1;
    wire   [0:0] icmp_ln133_87_fu_2937_p2;
    wire   [0:0] icmp_ln133_86_fu_2931_p2;
    wire   [10:0] tmp_233_fu_2917_p4;
    wire   [51:0] trunc_ln133_43_fu_2927_p1;
    wire   [0:0] icmp_ln133_89_fu_2955_p2;
    wire   [0:0] icmp_ln133_88_fu_2949_p2;
    wire   [0:0] or_ln133_43_fu_2961_p2;
    wire   [0:0] and_ln133_42_fu_2967_p2;
    wire   [0:0] and_ln133_43_fu_2973_p2;
    wire   [63:0] bitcast_ln135_42_fu_2985_p1;
    wire   [63:0] bitcast_ln135_43_fu_3003_p1;
    wire   [10:0] tmp_237_fu_2989_p4;
    wire   [51:0] trunc_ln135_42_fu_2999_p1;
    wire   [0:0] icmp_ln135_87_fu_3026_p2;
    wire   [0:0] icmp_ln135_86_fu_3020_p2;
    wire   [10:0] tmp_238_fu_3006_p4;
    wire   [51:0] trunc_ln135_43_fu_3016_p1;
    wire   [0:0] icmp_ln135_89_fu_3044_p2;
    wire   [0:0] icmp_ln135_88_fu_3038_p2;
    wire   [0:0] or_ln135_42_fu_3032_p2;
    wire   [0:0] or_ln135_43_fu_3050_p2;
    wire   [0:0] and_ln135_42_fu_3056_p2;
    wire   [0:0] and_ln135_43_fu_3062_p2;
    wire   [63:0] bitcast_ln136_17_fu_3075_p1;
    wire   [10:0] tmp_240_fu_3078_p4;
    wire   [51:0] trunc_ln136_17_fu_3088_p1;
    wire   [0:0] icmp_ln136_37_fu_3098_p2;
    wire   [0:0] icmp_ln136_36_fu_3092_p2;
    wire   [0:0] or_ln136_17_fu_3104_p2;
    wire   [0:0] and_ln136_39_fu_3110_p2;
    wire   [0:0] and_ln136_40_fu_3116_p2;
    wire   [63:0] bitcast_ln134_17_fu_3129_p1;
    wire   [10:0] tmp_235_fu_3132_p4;
    wire   [51:0] trunc_ln134_17_fu_3142_p1;
    wire   [0:0] icmp_ln134_37_fu_3152_p2;
    wire   [0:0] icmp_ln134_36_fu_3146_p2;
    wire   [0:0] or_ln134_17_fu_3158_p2;
    wire   [0:0] and_ln134_39_fu_3164_p2;
    wire   [0:0] and_ln134_40_fu_3169_p2;
    wire   [63:0] bitcast_ln135_44_fu_3181_p1;
    wire   [63:0] bitcast_ln135_45_fu_3198_p1;
    wire   [10:0] tmp_247_fu_3184_p4;
    wire   [51:0] trunc_ln135_44_fu_3194_p1;
    wire   [0:0] icmp_ln135_91_fu_3221_p2;
    wire   [0:0] icmp_ln135_90_fu_3215_p2;
    wire   [10:0] tmp_248_fu_3201_p4;
    wire   [51:0] trunc_ln135_45_fu_3211_p1;
    wire   [0:0] icmp_ln135_93_fu_3239_p2;
    wire   [0:0] icmp_ln135_92_fu_3233_p2;
    wire   [0:0] or_ln135_44_fu_3227_p2;
    wire   [0:0] or_ln135_45_fu_3245_p2;
    wire   [0:0] and_ln135_44_fu_3251_p2;
    wire   [0:0] and_ln135_45_fu_3257_p2;
    wire   [63:0] bitcast_ln136_18_fu_3269_p1;
    wire   [10:0] tmp_250_fu_3272_p4;
    wire   [51:0] trunc_ln136_18_fu_3282_p1;
    wire   [0:0] icmp_ln136_39_fu_3292_p2;
    wire   [0:0] icmp_ln136_38_fu_3286_p2;
    wire   [0:0] or_ln136_18_fu_3298_p2;
    wire   [0:0] and_ln136_41_fu_3304_p2;
    wire   [0:0] and_ln136_42_fu_3310_p2;
    wire   [63:0] bitcast_ln133_44_fu_3322_p1;
    wire   [63:0] bitcast_ln133_45_fu_3339_p1;
    wire   [10:0] tmp_242_fu_3325_p4;
    wire   [51:0] trunc_ln133_44_fu_3335_p1;
    wire   [0:0] icmp_ln133_91_fu_3362_p2;
    wire   [0:0] icmp_ln133_90_fu_3356_p2;
    wire   [10:0] tmp_243_fu_3342_p4;
    wire   [51:0] trunc_ln133_45_fu_3352_p1;
    wire   [0:0] icmp_ln133_93_fu_3380_p2;
    wire   [0:0] icmp_ln133_92_fu_3374_p2;
    wire   [0:0] or_ln133_44_fu_3368_p2;
    wire   [0:0] or_ln133_45_fu_3386_p2;
    wire   [0:0] and_ln133_44_fu_3392_p2;
    wire   [0:0] and_ln133_45_fu_3398_p2;
    wire   [63:0] bitcast_ln134_18_fu_3410_p1;
    wire   [10:0] tmp_245_fu_3413_p4;
    wire   [51:0] trunc_ln134_18_fu_3423_p1;
    wire   [0:0] icmp_ln134_39_fu_3433_p2;
    wire   [0:0] icmp_ln134_38_fu_3427_p2;
    wire   [0:0] or_ln134_18_fu_3439_p2;
    wire   [0:0] and_ln134_41_fu_3445_p2;
    wire   [0:0] and_ln134_42_fu_3451_p2;
    wire   [63:0] bitcast_ln139_fu_3463_p1;
    wire   [63:0] bitcast_ln139_5_fu_3480_p1;
    wire   [10:0] tmp_252_fu_3466_p4;
    wire   [51:0] trunc_ln139_fu_3476_p1;
    wire   [0:0] icmp_ln139_11_fu_3503_p2;
    wire   [0:0] icmp_ln139_fu_3497_p2;
    wire   [10:0] tmp_253_fu_3483_p4;
    wire   [51:0] trunc_ln139_5_fu_3493_p1;
    wire   [0:0] icmp_ln139_13_fu_3521_p2;
    wire   [0:0] icmp_ln139_12_fu_3515_p2;
    wire   [0:0] or_ln139_fu_3509_p2;
    wire   [0:0] or_ln139_5_fu_3527_p2;
    wire   [63:0] bitcast_ln139_6_fu_3539_p1;
    wire   [10:0] tmp_255_fu_3542_p4;
    wire   [51:0] trunc_ln139_6_fu_3552_p1;
    wire   [0:0] icmp_ln139_15_fu_3562_p2;
    wire   [0:0] icmp_ln139_14_fu_3556_p2;
    wire   [0:0] or_ln139_6_fu_3568_p2;
    wire   [0:0] and_ln139_11_fu_3574_p2;
    wire   [63:0] bitcast_ln140_fu_3585_p1;
    wire   [10:0] tmp_257_fu_3588_p4;
    wire   [51:0] trunc_ln140_fu_3598_p1;
    wire   [0:0] icmp_ln140_3_fu_3608_p2;
    wire   [0:0] icmp_ln140_fu_3602_p2;
    wire   [0:0] or_ln140_7_fu_3614_p2;
    wire   [0:0] and_ln140_9_fu_3620_p2;
    wire   [0:0] and_ln140_12_fu_3637_p2;
    wire   [0:0] and_ln141_fu_3642_p2;
    wire   [0:0] and_ln140_10_fu_3626_p2;
    wire   [0:0] or_ln140_fu_3647_p2;
    wire   [0:0] and_ln142_3_fu_3659_p2;
    wire   [0:0] and_ln142_fu_3664_p2;
    wire   [0:0] and_ln139_10_fu_3674_p2;
    wire   [0:0] and_ln139_fu_3678_p2;
    reg   [4:0] grp_fu_790_opcode;
    wire    ap_block_pp0_stage5_00001;
    wire    ap_block_pp0_stage6_00001;
    wire    ap_block_pp0_stage7_00001;
    wire    ap_block_pp0_stage8_00001;
    wire    ap_block_pp0_stage9_00001;
    wire    ap_block_pp0_stage10_00001;
    wire    ap_block_pp0_stage11_00001;
    wire    ap_block_pp0_stage12_00001;
    wire    ap_block_pp0_stage13_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage4_00001;
    reg   [4:0] grp_fu_794_opcode;
    reg   [4:0] grp_fu_798_opcode;
    reg   [13:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to4;
    wire    ap_block_pp0_stage1_subdone;
    reg    ap_idle_pp0_0to3;
    reg    ap_reset_idle_pp0;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_enable_pp0;
    wire   [6:0] mul_ln120_fu_984_p00;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 14'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
    end

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1246 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_746_p0),
        .din1(grp_fu_746_p1),
        .ce(1'b1),
        .dout(grp_fu_746_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1247 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_751_p0),
        .din1(grp_fu_751_p1),
        .ce(1'b1),
        .dout(grp_fu_751_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1248 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_756_p0),
        .din1(grp_fu_756_p1),
        .ce(1'b1),
        .dout(grp_fu_756_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1249 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_761_p0),
        .din1(grp_fu_761_p1),
        .ce(1'b1),
        .dout(grp_fu_761_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1250 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_766_p0),
        .din1(grp_fu_766_p1),
        .ce(1'b1),
        .dout(grp_fu_766_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1251 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_771_p0),
        .din1(grp_fu_771_p1),
        .ce(1'b1),
        .dout(grp_fu_771_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1252 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_776_p0),
        .din1(grp_fu_776_p1),
        .ce(1'b1),
        .dout(grp_fu_776_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1253 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_781_p0),
        .din1(grp_fu_781_p1),
        .ce(1'b1),
        .dout(grp_fu_781_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1254 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_790_p0),
        .din1(grp_fu_790_p1),
        .ce(1'b1),
        .opcode(grp_fu_790_opcode),
        .dout(grp_fu_790_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1255 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_794_p0),
        .din1(grp_fu_794_p1),
        .ce(1'b1),
        .opcode(grp_fu_794_opcode),
        .dout(grp_fu_794_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1256 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_798_p0),
        .din1(grp_fu_798_p1),
        .ce(1'b1),
        .opcode(grp_fu_798_opcode),
        .dout(grp_fu_798_p2)
    );

    main_mul_2ns_6ns_7_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(2),
        .din1_WIDTH(6),
        .dout_WIDTH(7)
    ) mul_2ns_6ns_7_1_1_U1257 (
        .din0(mul_ln120_fu_984_p0),
        .din1(mul_ln120_fu_984_p1),
        .dout(mul_ln120_fu_984_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                ap_enable_reg_pp0_iter4 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage9_11001) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                reg_807 <= p1_q0;
            end else if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                reg_807 <= p1_q1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage9_11001) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                reg_814 <= p1_q1;
            end else if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                reg_814 <= p1_q0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            and_ln133_reg_4557 <= and_ln133_fu_1327_p2;
            max2_reg_4568 <= max2_fu_1417_p3;
            min2_20_reg_4575 <= min2_20_fu_1431_p3;
            mul25_7_2_reg_4467_pp0_iter2_reg <= mul25_7_2_reg_4467;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            and_ln139_12_reg_4888 <= and_ln139_12_fu_3580_p2;
            and_ln139_9_reg_4883 <= and_ln139_9_fu_3533_p2;
            and_ln140_11_reg_4894 <= and_ln140_11_fu_3631_p2;
            and_ln140_reg_4899 <= and_ln140_fu_3653_p2;
            max1_29_reg_4721 <= max1_29_fu_2406_p3;
            max2_29_reg_4728 <= max2_29_fu_2496_p3;
            min2_24_reg_4735 <= min2_24_fu_2550_p3;
            mul_ln120_reg_3688 <= mul_ln120_fu_984_p2;
            or_ln133_38_reg_4716 <= or_ln133_38_fu_2370_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_port_reg_p_read  <= p_read;
            ap_port_reg_p_read1 <= p_read1;
            ap_port_reg_p_read2 <= p_read2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            max1_1_reg_4487 <= grp_fu_746_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            max1_26_reg_4614 <= max1_26_fu_1548_p3;
            max2_26_reg_4621 <= max2_26_fu_1638_p3;
            min2_21_reg_4628 <= min2_21_fu_1692_p3;
            or_ln133_32_reg_4609 <= or_ln133_32_fu_1512_p2;
            p_read_64_reg_4079 <= ap_port_reg_p_read2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            max1_27_reg_4647 <= max1_27_fu_1835_p3;
            max2_27_reg_4654 <= max2_27_fu_1925_p3;
            min2_22_reg_4661 <= min2_22_fu_1979_p3;
            or_ln133_34_reg_4642 <= or_ln133_34_fu_1799_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            max1_28_reg_4680 <= max1_28_fu_2121_p3;
            max2_28_reg_4687 <= max2_28_fu_2210_p3;
            min2_23_reg_4694 <= min2_23_fu_2264_p3;
            or_ln133_36_reg_4675 <= or_ln133_36_fu_2085_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            max1_30_reg_4772 <= max1_30_fu_2693_p3;
            max2_30_reg_4779 <= max2_30_fu_2783_p3;
            min2_25_reg_4786 <= min2_25_fu_2837_p3;
            or_ln133_40_reg_4767 <= or_ln133_40_fu_2657_p2;
            p_read83_reg_4003 <= ap_port_reg_p_read;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            max1_31_reg_4805 <= max1_31_fu_2979_p3;
            max2_31_reg_4812 <= max2_31_fu_3068_p3;
            min2_26_reg_4819 <= min2_26_fu_3122_p3;
            or_ln133_42_reg_4800 <= or_ln133_42_fu_2943_p2;
            p_read_65_reg_4031 <= ap_port_reg_p_read1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            max1_32_reg_4848 <= max1_32_fu_3404_p3;
            min1_21_reg_4635 <= min1_21_fu_1745_p3;
            min1_27_reg_4855 <= min1_27_fu_3457_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            max1_33_reg_4292 <= grp_fu_746_p2;
            mul20_8_reg_4302 <= grp_fu_771_p2;
            mul25_4_1_reg_4312 <= grp_fu_776_p2;
            mul25_7_reg_4317 <= grp_fu_781_p2;
            mul_2_reg_4297 <= grp_fu_766_p2;
            n2_3_reg_4307 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            max1_reg_4582 <= max1_fu_1443_p3;
            max2_32_reg_4833 <= max2_32_fu_3263_p3;
            min1_20_reg_4589 <= min1_20_fu_1457_p3;
            min2_27_reg_4841 <= min2_27_fu_3316_p3;
            mul20_7_2_reg_4482_pp0_iter2_reg <= mul20_7_2_reg_4482;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            min1_22_reg_4668 <= min1_22_fu_2032_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            min1_23_reg_4701 <= min1_23_fu_2317_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            min1_24_reg_4760 <= min1_24_fu_2603_p3;
            or_ln140_8_reg_4909 <= or_ln140_8_fu_3669_p2;
            p2_0_0_load_reg_3868 <= p2_0_0_q0;
            p2_0_1_load_reg_3873 <= p2_0_1_q0;
            p2_0_2_load_reg_3878 <= p2_0_2_q0;
            p2_1_0_load_reg_3883 <= p2_1_0_q0;
            p2_1_1_load_reg_3888 <= p2_1_1_q0;
            p2_1_2_load_reg_3893 <= p2_1_2_q0;
            p2_2_0_load_reg_3898 <= p2_2_0_q0;
            p2_2_1_load_reg_3903 <= p2_2_1_q0;
            p2_2_2_load_reg_3908 <= p2_2_2_q0;
            p2_3_0_load_reg_3913 <= p2_3_0_q0;
            p2_3_1_load_reg_3918 <= p2_3_1_q0;
            p2_3_2_load_reg_3923 <= p2_3_2_q0;
            p2_4_0_load_reg_3928 <= p2_4_0_q0;
            p2_4_1_load_reg_3933 <= p2_4_1_q0;
            p2_4_2_load_reg_3938 <= p2_4_2_q0;
            p2_5_0_load_reg_3943 <= p2_5_0_q0;
            p2_5_1_load_reg_3948 <= p2_5_1_q0;
            p2_5_2_load_reg_3953 <= p2_5_2_q0;
            p2_6_0_load_reg_3958 <= p2_6_0_q0;
            p2_6_1_load_reg_3963 <= p2_6_1_q0;
            p2_6_2_load_reg_3968 <= p2_6_2_q0;
            p2_7_0_load_reg_3973 <= p2_7_0_q0;
            p2_7_1_load_reg_3978 <= p2_7_1_q0;
            p2_7_2_load_reg_3983 <= p2_7_2_q0;
            p2_8_0_load_reg_3988 <= p2_8_0_q0;
            p2_8_1_load_reg_3993 <= p2_8_1_q0;
            p2_8_2_load_reg_3998 <= p2_8_2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            min1_25_reg_4793 <= min1_25_fu_2890_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            min1_26_reg_4826 <= min1_26_fu_3175_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            mul1_reg_4132 <= grp_fu_766_p2;
            mul20_1_reg_4137 <= grp_fu_771_p2;
            mul25_2_reg_4142 <= grp_fu_776_p2;
            mul25_3_reg_4147 <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            mul20_1_1_reg_4222 <= grp_fu_766_p2;
            mul20_4_reg_4232   <= grp_fu_776_p2;
            mul25_2_1_reg_4227 <= grp_fu_771_p2;
            mul25_5_reg_4237   <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            mul20_1_2_reg_4357 <= grp_fu_766_p2;
            mul20_5_1_reg_4377 <= grp_fu_776_p2;
            mul25_2_2_reg_4367 <= grp_fu_771_p2;
            mul25_6_1_reg_4382 <= grp_fu_781_p2;
            n1_6_reg_4362 <= grp_fu_746_p2;
            n1_9_reg_4372 <= grp_fu_751_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            mul20_2_1_reg_4252 <= grp_fu_766_p2;
            mul20_5_reg_4262   <= grp_fu_776_p2;
            mul25_3_1_reg_4257 <= grp_fu_771_p2;
            mul25_6_reg_4267   <= grp_fu_781_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul20_2_2_reg_4387 <= grp_fu_766_p2;
            mul20_6_1_reg_4402 <= grp_fu_776_p2;
            mul25_3_2_reg_4392 <= grp_fu_771_p2;
            mul25_7_1_reg_4407 <= grp_fu_781_p2;
            n2_40_reg_4397 <= grp_fu_746_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            mul20_2_reg_4172 <= grp_fu_776_p2;
            mul20_3_reg_4177 <= grp_fu_781_p2;
            mul25_s_reg_4167 <= grp_fu_771_p2;
            mul6_1_reg_4162  <= grp_fu_766_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            mul20_3_1_reg_4282 <= grp_fu_776_p2;
            mul20_6_reg_4287 <= grp_fu_781_p2;
            mul25_8_reg_4277 <= grp_fu_771_p2;
            mul6_2_reg_4272 <= grp_fu_766_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            mul20_3_2_reg_4412 <= grp_fu_766_p2;
            mul20_7_1_reg_4437 <= grp_fu_781_p2;
            mul25_4_2_reg_4422 <= grp_fu_771_p2;
            mul25_5_2_reg_4432 <= grp_fu_776_p2;
            n1_40_reg_4417 <= grp_fu_746_p2;
            n2_43_reg_4427 <= grp_fu_751_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            mul20_4_1_reg_4342 <= grp_fu_771_p2;
            mul20_7_reg_4352 <= grp_fu_781_p2;
            mul25_1_2_reg_4332 <= grp_fu_766_p2;
            mul25_5_1_reg_4347 <= grp_fu_776_p2;
            n1_3_reg_4327 <= grp_fu_751_p2;
            n1_reg_4322 <= grp_fu_746_p2;
            n2_6_reg_4337 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            mul20_4_2_reg_4442 <= grp_fu_766_p2;
            mul20_5_2_reg_4452 <= grp_fu_771_p2;
            mul25_6_2_reg_4462 <= grp_fu_776_p2;
            mul25_7_2_reg_4467 <= grp_fu_781_p2;
            n1_43_reg_4447 <= grp_fu_746_p2;
            n2_46_reg_4457 <= grp_fu_751_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            mul20_6_2_reg_4477 <= grp_fu_766_p2;
            mul20_7_2_reg_4482 <= grp_fu_771_p2;
            n1_46_reg_4472 <= grp_fu_746_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            mul20_s_reg_4197 <= grp_fu_771_p2;
            mul25_1_1_reg_4202 <= grp_fu_776_p2;
            mul25_4_reg_4207 <= grp_fu_781_p2;
            mul_1_reg_4192 <= grp_fu_766_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            mul25_1_reg_4117 <= grp_fu_781_p2;
            mul2_reg_4107 <= grp_fu_776_p2;
            mul6_reg_4102 <= grp_fu_771_p2;
            mul_reg_4097 <= grp_fu_766_p2;
            p1_load_5_reg_4112 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            n1_1_reg_4492  <= grp_fu_746_p2;
            n1_4_reg_4497  <= grp_fu_751_p2;
            n2_38_reg_4502 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            n1_38_reg_4512 <= grp_fu_751_p2;
            n1_49_reg_4517 <= grp_fu_756_p2;
            n1_7_reg_4507  <= grp_fu_746_p2;
            n2_49_reg_4522 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            n1_39_reg_4596 <= grp_fu_751_p2;
            n2_50_reg_4604 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            n1_41_reg_4532 <= grp_fu_746_p2;
            n2_44_reg_4537 <= grp_fu_751_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            n1_44_reg_4542 <= grp_fu_746_p2;
            n2_47_reg_4547 <= grp_fu_751_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            n1_47_reg_4552 <= grp_fu_746_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            n1_48_reg_4708 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            n1_51_reg_4742 <= grp_fu_751_p2;
            n2_51_reg_4751 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            n2_41_reg_4527 <= grp_fu_746_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            reg_802 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_821 <= p1_q0;
            reg_827 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_833 <= p1_q0;
            reg_838 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            reg_844 <= p1_q0;
            reg_849 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_855 <= p1_q0;
            reg_860 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_866 <= p1_q0;
            reg_872 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            reg_878 <= grp_fu_751_p2;
            reg_884 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            reg_891 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_898 <= grp_fu_751_p2;
            reg_904 <= grp_fu_756_p2;
            reg_911 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)))) begin
            reg_918 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_924 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_930 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            reg_938 <= grp_fu_761_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            reg_944 <= grp_fu_756_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            tmp_176_reg_4563 <= grp_fu_790_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            tmp_254_reg_4904 <= grp_fu_794_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            tmp_256_reg_4863 <= grp_fu_794_p2;
            tmp_258_reg_4868 <= grp_fu_798_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            tmp_259_reg_4873 <= grp_fu_794_p2;
            tmp_260_reg_4878 <= grp_fu_798_p2;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to3 = 1'b1;
        end else begin
            ap_idle_pp0_0to3 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to4 = 1'b1;
        end else begin
            ap_idle_pp0_1to4 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0_0to3 == 1'b1) & (ap_start == 1'b0))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_746_p0 = n1_46_reg_4472;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_746_p0 = n1_43_reg_4447;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_746_p0 = n1_40_reg_4417;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_746_p0 = n2_40_reg_4397;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_746_p0 = n1_6_reg_4362;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_746_p0 = n1_reg_4322;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_746_p0 = max1_33_reg_4292;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_746_p0 = mul20_6_reg_4287;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_746_p0 = mul20_5_reg_4262;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_746_p0 = mul20_4_reg_4232;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_746_p0 = mul25_4_reg_4207;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_746_p0 = mul20_2_reg_4172;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_746_p0 = mul1_reg_4132;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_746_p0 = mul_reg_4097;
        end else begin
            grp_fu_746_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_746_p1 = mul20_6_1_reg_4402;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_746_p1 = mul20_5_1_reg_4377;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_746_p1 = mul20_4_1_reg_4342;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_746_p1 = mul25_4_1_reg_4312;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_746_p1 = mul20_2_1_reg_4252;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_746_p1 = mul20_s_reg_4197;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_746_p1 = mul_1_reg_4192;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_746_p1 = 64'd0;
        end else begin
            grp_fu_746_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_751_p0 = reg_924;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_751_p0 = n1_41_reg_4532;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_751_p0 = n1_38_reg_4512;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_751_p0 = n1_1_reg_4492;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_751_p0 = n2_46_reg_4457;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_751_p0 = n2_43_reg_4427;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_751_p0 = n1_9_reg_4372;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_751_p0 = n1_3_reg_4327;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_751_p0 = reg_878;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_751_p0 = mul25_6_reg_4267;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_751_p0 = mul25_5_reg_4237;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_751_p0 = mul20_3_reg_4177;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_751_p0 = mul20_1_reg_4137;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_751_p0 = mul6_reg_4102;
        end else begin
            grp_fu_751_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_751_p1 = mul20_7_2_reg_4482_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_751_p1 = mul20_4_2_reg_4442;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_751_p1 = mul20_3_2_reg_4412;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_751_p1 = mul20_8_reg_4302;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_751_p1 = mul25_6_1_reg_4382;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_751_p1 = mul25_5_1_reg_4347;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_751_p1 = mul20_3_1_reg_4282;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_751_p1 = mul20_1_1_reg_4222;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_751_p1 = mul6_1_reg_4162;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_751_p1 = 64'd0;
        end else begin
            grp_fu_751_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_756_p0 = n2_50_reg_4604;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_756_p0 = n1_47_reg_4552;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_756_p0 = n1_44_reg_4542;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_756_p0 = n2_41_reg_4527;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_756_p0 = n1_49_reg_4517;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_756_p0 = n1_7_reg_4507;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_756_p0 = n1_4_reg_4497;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_756_p0 = reg_904;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_756_p0 = max1_1_reg_4487;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_756_p0 = mul20_7_reg_4352;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_756_p0 = n2_6_reg_4337;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_756_p0 = reg_884;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_756_p0 = mul25_2_reg_4142;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_756_p0 = mul2_reg_4107;
        end else begin
            grp_fu_756_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_756_p1 = mul25_7_2_reg_4467_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_756_p1 = mul20_6_2_reg_4477;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_756_p1 = mul20_5_2_reg_4452;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_756_p1 = mul25_4_2_reg_4422;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_756_p1 = mul20_7_1_reg_4437;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_756_p1 = mul20_2_2_reg_4387;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_756_p1 = mul20_1_2_reg_4357;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_756_p1 = mul25_8_reg_4277;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_756_p1 = mul_2_reg_4297;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_756_p1 = mul25_2_1_reg_4227;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_756_p1 = mul25_s_reg_4167;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_756_p1 = 64'd0;
        end else begin
            grp_fu_756_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_761_p0 = n2_47_reg_4547;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_761_p0 = n2_44_reg_4537;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_761_p0 = n2_49_reg_4522;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_761_p0 = n2_38_reg_4502;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_761_p0 = reg_918;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_761_p0 = reg_911;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_761_p0 = reg_898;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_761_p0 = mul25_7_reg_4317;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_761_p0 = reg_891;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_761_p0 = n2_3_reg_4307;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_761_p0 = mul25_3_reg_4147;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_761_p0 = mul25_1_reg_4117;
        end else begin
            grp_fu_761_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_761_p1 = mul25_6_2_reg_4462;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_761_p1 = mul25_5_2_reg_4432;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_761_p1 = mul25_7_1_reg_4407;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_761_p1 = mul25_3_2_reg_4392;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_761_p1 = mul25_2_2_reg_4367;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_761_p1 = mul25_1_2_reg_4332;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_761_p1 = mul6_2_reg_4272;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_761_p1 = mul25_3_1_reg_4257;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_761_p1 = mul25_1_1_reg_4202;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_761_p1 = 64'd0;
        end else begin
            grp_fu_761_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_766_p0 = reg_866;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_766_p0 = reg_821;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_766_p0 = p2_2_2_load_reg_3908;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_766_p0 = p2_0_2_load_reg_3878;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_766_p0 = reg_855;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_766_p0 = reg_844;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_766_p0 = reg_833;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_766_p0 = p2_0_1_load_reg_3873;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_766_p0 = reg_807;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_766_p0 = reg_802;
        end else begin
            grp_fu_766_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_766_p1 = p_read_64_reg_4079;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_766_p1 = ap_port_reg_p_read2;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_766_p1 = p_read_65_reg_4031;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_766_p1 = ap_port_reg_p_read1;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_766_p1 = p_read83_reg_4003;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_766_p1 = ap_port_reg_p_read;
        end else begin
            grp_fu_766_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_771_p0 = reg_872;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_771_p0 = reg_860;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_771_p0 = p2_5_2_load_reg_3953;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_771_p0 = p2_4_2_load_reg_3938;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_771_p0 = p2_3_2_load_reg_3923;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_771_p0 = reg_807;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_771_p0 = p1_load_5_reg_4112;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_771_p0 = p2_1_2_load_reg_3893;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_771_p0 = p2_4_1_load_reg_3933;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_771_p0 = p2_3_1_load_reg_3918;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_771_p0 = reg_838;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_771_p0 = p2_1_1_load_reg_3888;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_771_p0 = reg_814;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_771_p0 = p2_0_0_load_reg_3868;
        end else begin
            grp_fu_771_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_771_p1 = p_read_64_reg_4079;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_771_p1 = ap_port_reg_p_read2;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_771_p1 = p_read_65_reg_4031;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_771_p1 = ap_port_reg_p_read1;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_771_p1 = p_read83_reg_4003;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_771_p1 = ap_port_reg_p_read;
        end else begin
            grp_fu_771_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_776_p0 = p2_7_2_load_reg_3983;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_776_p0 = p2_6_2_load_reg_3968;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_776_p0 = reg_838;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_776_p0 = reg_827;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_776_p0 = p2_6_1_load_reg_3963;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_776_p0 = p2_5_1_load_reg_3948;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_776_p0 = reg_866;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_776_p0 = reg_860;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_776_p0 = reg_849;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_776_p0 = p2_2_1_load_reg_3903;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_776_p0 = reg_821;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_776_p0 = p2_3_0_load_reg_3913;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_776_p0 = p2_1_0_load_reg_3883;
        end else begin
            grp_fu_776_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_776_p1 = p_read_64_reg_4079;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_776_p1 = p_read_65_reg_4031;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_776_p1 = p_read83_reg_4003;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_776_p1 = ap_port_reg_p_read;
        end else begin
            grp_fu_776_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_781_p0 = p2_8_2_load_reg_3998;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_781_p0 = reg_849;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_781_p0 = p2_8_1_load_reg_3993;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_781_p0 = p2_7_1_load_reg_3978;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_781_p0 = reg_814;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_781_p0 = p2_8_0_load_reg_3988;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_781_p0 = reg_872;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_781_p0 = p2_7_0_load_reg_3973;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_781_p0 = p2_6_0_load_reg_3958;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_781_p0 = p2_5_0_load_reg_3943;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_781_p0 = reg_827;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_781_p0 = p2_4_0_load_reg_3928;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_781_p0 = p2_2_0_load_reg_3898;
        end else begin
            grp_fu_781_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_781_p1 = p_read_64_reg_4079;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_781_p1 = p_read_65_reg_4031;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_781_p1 = p_read83_reg_4003;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_781_p1 = ap_port_reg_p_read;
        end else begin
            grp_fu_781_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_790_opcode = 5'd4;
        end else if ((((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_790_opcode = 5'd2;
        end else begin
            grp_fu_790_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_790_p0 = n1_48_reg_4708;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_790_p0 = reg_878;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_790_p0 = n1_39_reg_4596;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_790_p0 = reg_944;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_790_p0 = reg_918;
        end else if ((((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_790_p0 = reg_898;
        end else begin
            grp_fu_790_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_790_p1 = min1_25_reg_4793;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_790_p1 = max1_30_reg_4772;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_790_p1 = min1_24_reg_4760;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_790_p1 = max1_29_reg_4721;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_790_p1 = min1_23_reg_4701;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_790_p1 = max1_28_reg_4680;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_790_p1 = min1_22_reg_4668;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_790_p1 = max1_27_reg_4647;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_790_p1 = min1_21_reg_4635;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_790_p1 = max1_26_reg_4614;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_790_p1 = min1_20_reg_4589;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_790_p1 = max1_fu_1443_p3;
        end else if ((((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_790_p1 = reg_924;
        end else begin
            grp_fu_790_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_794_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_794_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_794_opcode = 5'd2;
        end else begin
            grp_fu_794_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_794_p0 = min1_27_reg_4855;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_794_p0 = max1_32_reg_4848;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_794_p0 = n1_51_reg_4742;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_794_p0 = n2_51_reg_4751;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_794_p0 = reg_891;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_794_p0 = reg_884;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_794_p0 = reg_930;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_794_p0 = reg_938;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_794_p0 = reg_911;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_794_p0 = reg_904;
        end else begin
            grp_fu_794_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_794_p1 = max2_32_reg_4833;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_794_p1 = min2_27_reg_4841;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_794_p1 = max1_31_reg_4805;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_794_p1 = max2_31_reg_4812;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_794_p1 = max2_30_reg_4779;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_794_p1 = max2_29_reg_4728;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_794_p1 = max2_28_reg_4687;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_794_p1 = max2_27_reg_4654;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_794_p1 = max2_26_reg_4621;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_794_p1 = max2_reg_4568;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_794_p1 = reg_930;
        end else begin
            grp_fu_794_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_798_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_798_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_798_opcode = 5'd4;
        end else begin
            grp_fu_798_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_798_p0 = min2_27_reg_4841;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_798_p0 = max2_32_reg_4833;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_798_p0 = min1_27_reg_4855;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_798_p0 = n1_51_reg_4742;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_798_p0 = n2_51_reg_4751;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_798_p0 = reg_891;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_798_p0 = reg_884;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_798_p0 = reg_930;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_798_p0 = reg_938;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_798_p0 = reg_911;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_798_p0 = reg_904;
        end else begin
            grp_fu_798_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_798_p1 = min1_27_reg_4855;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_798_p1 = max1_32_reg_4848;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_798_p1 = max2_32_reg_4833;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_798_p1 = min1_26_reg_4826;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_798_p1 = min2_26_reg_4819;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_798_p1 = min2_25_reg_4786;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_798_p1 = min2_24_reg_4735;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_798_p1 = min2_23_reg_4694;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_798_p1 = min2_22_reg_4661;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_798_p1 = min2_21_reg_4628;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_798_p1 = min2_20_reg_4575;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_798_p1 = reg_930;
        end else begin
            grp_fu_798_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address0 = zext_ln129_66_fu_1240_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address0 = zext_ln129_60_fu_1220_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address0 = zext_ln129_57_fu_1200_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address0 = zext_ln129_54_fu_1180_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address0 = zext_ln129_51_fu_1160_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address0 = zext_ln129_59_fu_1140_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address0 = zext_ln120_19_fu_1120_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address0 = zext_ln129_56_fu_1100_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address0 = zext_ln129_53_fu_1080_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address0 = zext_ln129_50_fu_1060_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address0 = zext_ln120_18_fu_1040_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address0 = zext_ln129_52_fu_1020_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address0 = zext_ln129_49_fu_1010_p1;
            end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                p1_address0 = zext_ln120_17_fu_990_p1;
            end else begin
                p1_address0 = 'bx;
            end
        end else begin
            p1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address1 = zext_ln129_69_fu_1250_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address1 = zext_ln129_63_fu_1230_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address1 = zext_ln129_68_fu_1210_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address1 = zext_ln129_65_fu_1190_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address1 = zext_ln129_62_fu_1170_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address1 = zext_ln129_67_fu_1150_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address1 = zext_ln129_48_fu_1130_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address1 = zext_ln129_64_fu_1110_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address1 = zext_ln129_61_fu_1090_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address1 = zext_ln129_58_fu_1070_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address1 = zext_ln129_47_fu_1050_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address1 = zext_ln129_55_fu_1030_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address1 = zext_ln129_fu_1000_p1;
            end else begin
                p1_address1 = 'bx;
            end
        end else begin
            p1_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            p1_ce0 = 1'b1;
        end else begin
            p1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            p1_ce1 = 1'b1;
        end else begin
            p1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_0_ce0 = 1'b1;
        end else begin
            p2_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_1_ce0 = 1'b1;
        end else begin
            p2_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_2_ce0 = 1'b1;
        end else begin
            p2_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_0_ce0 = 1'b1;
        end else begin
            p2_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_1_ce0 = 1'b1;
        end else begin
            p2_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_2_ce0 = 1'b1;
        end else begin
            p2_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_0_ce0 = 1'b1;
        end else begin
            p2_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_1_ce0 = 1'b1;
        end else begin
            p2_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_2_ce0 = 1'b1;
        end else begin
            p2_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_0_ce0 = 1'b1;
        end else begin
            p2_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_1_ce0 = 1'b1;
        end else begin
            p2_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_2_ce0 = 1'b1;
        end else begin
            p2_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_0_ce0 = 1'b1;
        end else begin
            p2_4_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_1_ce0 = 1'b1;
        end else begin
            p2_4_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_2_ce0 = 1'b1;
        end else begin
            p2_4_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_0_ce0 = 1'b1;
        end else begin
            p2_5_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_1_ce0 = 1'b1;
        end else begin
            p2_5_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_2_ce0 = 1'b1;
        end else begin
            p2_5_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_0_ce0 = 1'b1;
        end else begin
            p2_6_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_1_ce0 = 1'b1;
        end else begin
            p2_6_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_2_ce0 = 1'b1;
        end else begin
            p2_6_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_0_ce0 = 1'b1;
        end else begin
            p2_7_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_1_ce0 = 1'b1;
        end else begin
            p2_7_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_2_ce0 = 1'b1;
        end else begin
            p2_7_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_0_ce0 = 1'b1;
        end else begin
            p2_8_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_1_ce0 = 1'b1;
        end else begin
            p2_8_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_2_ce0 = 1'b1;
        end else begin
            p2_8_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_idle_pp0_1to4 == 1'b1) & (ap_start == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if (((1'b0 == ap_block_pp0_stage2_subdone) & (ap_reset_idle_pp0 == 1'b0))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else if (((1'b0 == ap_block_pp0_stage2_subdone) & (ap_reset_idle_pp0 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln120_9_fu_1115_p2 = (mul_ln120_reg_3688 + 7'd2);

    assign add_ln120_fu_1035_p2 = (mul_ln120_reg_3688 + 7'd1);

    assign add_ln129_47_fu_1045_p2 = (mul_ln120_reg_3688 + 7'd4);

    assign add_ln129_48_fu_1125_p2 = (mul_ln120_reg_3688 + 7'd5);

    assign add_ln129_49_fu_1005_p2 = (mul_ln120_reg_3688 + 7'd6);

    assign add_ln129_50_fu_1055_p2 = (mul_ln120_reg_3688 + 7'd7);

    assign add_ln129_51_fu_1155_p2 = (mul_ln120_reg_3688 + 7'd8);

    assign add_ln129_52_fu_1015_p2 = (mul_ln120_reg_3688 + 7'd9);

    assign add_ln129_53_fu_1075_p2 = (mul_ln120_reg_3688 + 7'd10);

    assign add_ln129_54_fu_1175_p2 = (mul_ln120_reg_3688 + 7'd11);

    assign add_ln129_55_fu_1025_p2 = (mul_ln120_reg_3688 + 7'd12);

    assign add_ln129_56_fu_1095_p2 = (mul_ln120_reg_3688 + 7'd13);

    assign add_ln129_57_fu_1195_p2 = (mul_ln120_reg_3688 + 7'd14);

    assign add_ln129_58_fu_1065_p2 = (mul_ln120_reg_3688 + 7'd15);

    assign add_ln129_59_fu_1135_p2 = (mul_ln120_reg_3688 + 7'd16);

    assign add_ln129_60_fu_1215_p2 = (mul_ln120_reg_3688 + 7'd17);

    assign add_ln129_61_fu_1085_p2 = (mul_ln120_reg_3688 + 7'd18);

    assign add_ln129_62_fu_1165_p2 = (mul_ln120_reg_3688 + 7'd19);

    assign add_ln129_63_fu_1225_p2 = (mul_ln120_reg_3688 + 7'd20);

    assign add_ln129_64_fu_1105_p2 = (mul_ln120_reg_3688 + 7'd21);

    assign add_ln129_65_fu_1185_p2 = (mul_ln120_reg_3688 + 7'd22);

    assign add_ln129_66_fu_1235_p2 = (mul_ln120_reg_3688 + 7'd23);

    assign add_ln129_67_fu_1145_p2 = (mul_ln120_reg_3688 + 7'd24);

    assign add_ln129_68_fu_1205_p2 = (mul_ln120_reg_3688 + 7'd25);

    assign add_ln129_69_fu_1245_p2 = (mul_ln120_reg_3688 + 7'd26);

    assign add_ln129_fu_995_p2 = (mul_ln120_reg_3688 + 7'd3);

    assign and_ln133_31_fu_1439_p2 = (tmp_176_reg_4563 & and_ln133_reg_4557);

    assign and_ln133_32_fu_1536_p2 = (or_ln133_33_fu_1530_p2 & or_ln133_32_fu_1512_p2);

    assign and_ln133_33_fu_1542_p2 = (grp_fu_790_p2 & and_ln133_32_fu_1536_p2);

    assign and_ln133_34_fu_1823_p2 = (or_ln133_35_fu_1817_p2 & or_ln133_34_fu_1799_p2);

    assign and_ln133_35_fu_1829_p2 = (grp_fu_790_p2 & and_ln133_34_fu_1823_p2);

    assign and_ln133_36_fu_2109_p2 = (or_ln133_37_fu_2103_p2 & or_ln133_36_fu_2085_p2);

    assign and_ln133_37_fu_2115_p2 = (grp_fu_790_p2 & and_ln133_36_fu_2109_p2);

    assign and_ln133_38_fu_2394_p2 = (or_ln133_39_fu_2388_p2 & or_ln133_38_fu_2370_p2);

    assign and_ln133_39_fu_2400_p2 = (grp_fu_790_p2 & and_ln133_38_fu_2394_p2);

    assign and_ln133_40_fu_2681_p2 = (or_ln133_41_fu_2675_p2 & or_ln133_40_fu_2657_p2);

    assign and_ln133_41_fu_2687_p2 = (grp_fu_790_p2 & and_ln133_40_fu_2681_p2);

    assign and_ln133_42_fu_2967_p2 = (or_ln133_43_fu_2961_p2 & or_ln133_42_fu_2943_p2);

    assign and_ln133_43_fu_2973_p2 = (grp_fu_790_p2 & and_ln133_42_fu_2967_p2);

    assign and_ln133_44_fu_3392_p2 = (or_ln133_45_fu_3386_p2 & or_ln133_44_fu_3368_p2);

    assign and_ln133_45_fu_3398_p2 = (grp_fu_794_p2 & and_ln133_44_fu_3392_p2);

    assign and_ln133_fu_1327_p2 = (or_ln133_fu_1303_p2 & or_ln133_31_fu_1321_p2);

    assign and_ln134_29_fu_1734_p2 = (or_ln134_fu_1728_p2 & or_ln133_32_reg_4609);

    assign and_ln134_30_fu_1739_p2 = (grp_fu_790_p2 & and_ln134_29_fu_1734_p2);

    assign and_ln134_31_fu_2021_p2 = (or_ln134_13_fu_2015_p2 & or_ln133_34_reg_4642);

    assign and_ln134_32_fu_2026_p2 = (grp_fu_790_p2 & and_ln134_31_fu_2021_p2);

    assign and_ln134_33_fu_2306_p2 = (or_ln134_14_fu_2300_p2 & or_ln133_36_reg_4675);

    assign and_ln134_34_fu_2311_p2 = (grp_fu_790_p2 & and_ln134_33_fu_2306_p2);

    assign and_ln134_35_fu_2592_p2 = (or_ln134_15_fu_2586_p2 & or_ln133_38_reg_4716);

    assign and_ln134_36_fu_2597_p2 = (grp_fu_790_p2 & and_ln134_35_fu_2592_p2);

    assign and_ln134_37_fu_2879_p2 = (or_ln134_16_fu_2873_p2 & or_ln133_40_reg_4767);

    assign and_ln134_38_fu_2884_p2 = (grp_fu_790_p2 & and_ln134_37_fu_2879_p2);

    assign and_ln134_39_fu_3164_p2 = (or_ln134_17_fu_3158_p2 & or_ln133_42_reg_4800);

    assign and_ln134_40_fu_3169_p2 = (grp_fu_790_p2 & and_ln134_39_fu_3164_p2);

    assign and_ln134_41_fu_3445_p2 = (or_ln134_18_fu_3439_p2 & or_ln133_44_fu_3368_p2);

    assign and_ln134_42_fu_3451_p2 = (grp_fu_798_p2 & and_ln134_41_fu_3445_p2);

    assign and_ln134_fu_1452_p2 = (grp_fu_790_p2 & and_ln133_reg_4557);

    assign and_ln135_31_fu_1411_p2 = (grp_fu_794_p2 & and_ln135_fu_1405_p2);

    assign and_ln135_32_fu_1626_p2 = (or_ln135_33_fu_1620_p2 & or_ln135_32_fu_1602_p2);

    assign and_ln135_33_fu_1632_p2 = (grp_fu_794_p2 & and_ln135_32_fu_1626_p2);

    assign and_ln135_34_fu_1913_p2 = (or_ln135_35_fu_1907_p2 & or_ln135_34_fu_1889_p2);

    assign and_ln135_35_fu_1919_p2 = (grp_fu_794_p2 & and_ln135_34_fu_1913_p2);

    assign and_ln135_36_fu_2198_p2 = (or_ln135_37_fu_2192_p2 & or_ln135_36_fu_2174_p2);

    assign and_ln135_37_fu_2204_p2 = (grp_fu_794_p2 & and_ln135_36_fu_2198_p2);

    assign and_ln135_38_fu_2484_p2 = (or_ln135_39_fu_2478_p2 & or_ln135_38_fu_2460_p2);

    assign and_ln135_39_fu_2490_p2 = (grp_fu_794_p2 & and_ln135_38_fu_2484_p2);

    assign and_ln135_40_fu_2771_p2 = (or_ln135_41_fu_2765_p2 & or_ln135_40_fu_2747_p2);

    assign and_ln135_41_fu_2777_p2 = (grp_fu_794_p2 & and_ln135_40_fu_2771_p2);

    assign and_ln135_42_fu_3056_p2 = (or_ln135_43_fu_3050_p2 & or_ln135_42_fu_3032_p2);

    assign and_ln135_43_fu_3062_p2 = (grp_fu_794_p2 & and_ln135_42_fu_3056_p2);

    assign and_ln135_44_fu_3251_p2 = (or_ln135_45_fu_3245_p2 & or_ln135_44_fu_3227_p2);

    assign and_ln135_45_fu_3257_p2 = (grp_fu_794_p2 & and_ln135_44_fu_3251_p2);

    assign and_ln135_fu_1405_p2 = (or_ln135_fu_1381_p2 & or_ln135_31_fu_1399_p2);

    assign and_ln136_29_fu_1680_p2 = (or_ln136_fu_1674_p2 & or_ln135_32_fu_1602_p2);

    assign and_ln136_30_fu_1686_p2 = (grp_fu_798_p2 & and_ln136_29_fu_1680_p2);

    assign and_ln136_31_fu_1967_p2 = (or_ln136_13_fu_1961_p2 & or_ln135_34_fu_1889_p2);

    assign and_ln136_32_fu_1973_p2 = (grp_fu_798_p2 & and_ln136_31_fu_1967_p2);

    assign and_ln136_33_fu_2252_p2 = (or_ln136_14_fu_2246_p2 & or_ln135_36_fu_2174_p2);

    assign and_ln136_34_fu_2258_p2 = (grp_fu_798_p2 & and_ln136_33_fu_2252_p2);

    assign and_ln136_35_fu_2538_p2 = (or_ln136_15_fu_2532_p2 & or_ln135_38_fu_2460_p2);

    assign and_ln136_36_fu_2544_p2 = (grp_fu_798_p2 & and_ln136_35_fu_2538_p2);

    assign and_ln136_37_fu_2825_p2 = (or_ln136_16_fu_2819_p2 & or_ln135_40_fu_2747_p2);

    assign and_ln136_38_fu_2831_p2 = (grp_fu_798_p2 & and_ln136_37_fu_2825_p2);

    assign and_ln136_39_fu_3110_p2 = (or_ln136_17_fu_3104_p2 & or_ln135_42_fu_3032_p2);

    assign and_ln136_40_fu_3116_p2 = (grp_fu_798_p2 & and_ln136_39_fu_3110_p2);

    assign and_ln136_41_fu_3304_p2 = (or_ln136_18_fu_3298_p2 & or_ln135_44_fu_3227_p2);

    assign and_ln136_42_fu_3310_p2 = (grp_fu_798_p2 & and_ln136_41_fu_3304_p2);

    assign and_ln136_fu_1425_p2 = (grp_fu_798_p2 & and_ln135_fu_1405_p2);

    assign and_ln139_10_fu_3674_p2 = (tmp_254_reg_4904 & and_ln139_9_reg_4883);

    assign and_ln139_11_fu_3574_p2 = (or_ln139_fu_3509_p2 & or_ln139_6_fu_3568_p2);

    assign and_ln139_12_fu_3580_p2 = (tmp_256_reg_4863 & and_ln139_11_fu_3574_p2);

    assign and_ln139_9_fu_3533_p2 = (or_ln139_fu_3509_p2 & or_ln139_5_fu_3527_p2);

    assign and_ln139_fu_3678_p2 = (and_ln139_12_reg_4888 & and_ln139_10_fu_3674_p2);

    assign and_ln140_10_fu_3626_p2 = (tmp_258_reg_4868 & and_ln140_9_fu_3620_p2);

    assign and_ln140_11_fu_3631_p2 = (or_ln140_7_fu_3614_p2 & or_ln139_6_fu_3568_p2);

    assign and_ln140_12_fu_3637_p2 = (tmp_259_reg_4873 & and_ln140_11_fu_3631_p2);

    assign and_ln140_9_fu_3620_p2 = (or_ln140_7_fu_3614_p2 & or_ln139_5_fu_3527_p2);

    assign and_ln140_fu_3653_p2 = (or_ln140_fu_3647_p2 & and_ln140_10_fu_3626_p2);

    assign and_ln141_fu_3642_p2 = (tmp_260_reg_4878 & and_ln139_9_fu_3533_p2);

    assign and_ln142_3_fu_3659_p2 = (grp_fu_798_p2 & and_ln140_11_reg_4894);

    assign and_ln142_fu_3664_p2 = (and_ln142_3_fu_3659_p2 & and_ln139_12_reg_4888);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_return = (or_ln140_8_reg_4909 | and_ln139_fu_3678_p2);

    assign bitcast_ln133_31_fu_1273_p1 = reg_924;

    assign bitcast_ln133_32_fu_1465_p1 = reg_918;

    assign bitcast_ln133_33_fu_1483_p1 = max1_reg_4582;

    assign bitcast_ln133_34_fu_1752_p1 = reg_944;

    assign bitcast_ln133_35_fu_1770_p1 = max1_26_reg_4614;

    assign bitcast_ln133_36_fu_2039_p1 = n1_39_reg_4596;

    assign bitcast_ln133_37_fu_2056_p1 = max1_27_reg_4647;

    assign bitcast_ln133_38_fu_2323_p1 = reg_878;

    assign bitcast_ln133_39_fu_2341_p1 = max1_28_reg_4680;

    assign bitcast_ln133_40_fu_2610_p1 = reg_944;

    assign bitcast_ln133_41_fu_2628_p1 = max1_29_reg_4721;

    assign bitcast_ln133_42_fu_2897_p1 = n1_48_reg_4708;

    assign bitcast_ln133_43_fu_2914_p1 = max1_30_reg_4772;

    assign bitcast_ln133_44_fu_3322_p1 = n1_51_reg_4742;

    assign bitcast_ln133_45_fu_3339_p1 = max1_31_reg_4805;

    assign bitcast_ln133_fu_1255_p1 = reg_898;

    assign bitcast_ln134_13_fu_1986_p1 = min1_21_reg_4635;

    assign bitcast_ln134_14_fu_2271_p1 = min1_22_reg_4668;

    assign bitcast_ln134_15_fu_2557_p1 = min1_23_reg_4701;

    assign bitcast_ln134_16_fu_2844_p1 = min1_24_reg_4760;

    assign bitcast_ln134_17_fu_3129_p1 = min1_25_reg_4793;

    assign bitcast_ln134_18_fu_3410_p1 = min1_26_reg_4826;

    assign bitcast_ln134_fu_1699_p1 = min1_20_reg_4589;

    assign bitcast_ln135_31_fu_1351_p1 = reg_930;

    assign bitcast_ln135_32_fu_1555_p1 = reg_911;

    assign bitcast_ln135_33_fu_1573_p1 = max2_reg_4568;

    assign bitcast_ln135_34_fu_1842_p1 = reg_938;

    assign bitcast_ln135_35_fu_1860_p1 = max2_26_reg_4621;

    assign bitcast_ln135_36_fu_2127_p1 = reg_930;

    assign bitcast_ln135_37_fu_2145_p1 = max2_27_reg_4654;

    assign bitcast_ln135_38_fu_2413_p1 = reg_884;

    assign bitcast_ln135_39_fu_2431_p1 = max2_28_reg_4687;

    assign bitcast_ln135_40_fu_2700_p1 = reg_891;

    assign bitcast_ln135_41_fu_2718_p1 = max2_29_reg_4728;

    assign bitcast_ln135_42_fu_2985_p1 = reg_938;

    assign bitcast_ln135_43_fu_3003_p1 = max2_30_reg_4779;

    assign bitcast_ln135_44_fu_3181_p1 = n2_51_reg_4751;

    assign bitcast_ln135_45_fu_3198_p1 = max2_31_reg_4812;

    assign bitcast_ln135_fu_1333_p1 = reg_904;

    assign bitcast_ln136_13_fu_1932_p1 = min2_21_reg_4628;

    assign bitcast_ln136_14_fu_2217_p1 = min2_22_reg_4661;

    assign bitcast_ln136_15_fu_2503_p1 = min2_23_reg_4694;

    assign bitcast_ln136_16_fu_2790_p1 = min2_24_reg_4735;

    assign bitcast_ln136_17_fu_3075_p1 = min2_25_reg_4786;

    assign bitcast_ln136_18_fu_3269_p1 = min2_26_reg_4819;

    assign bitcast_ln136_fu_1645_p1 = min2_20_reg_4575;

    assign bitcast_ln139_5_fu_3480_p1 = max2_32_reg_4833;

    assign bitcast_ln139_6_fu_3539_p1 = min2_27_reg_4841;

    assign bitcast_ln139_fu_3463_p1 = max1_32_reg_4848;

    assign bitcast_ln140_fu_3585_p1 = min1_27_reg_4855;

    assign icmp_ln133_63_fu_1297_p2 = ((trunc_ln133_fu_1269_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_64_fu_1309_p2 = ((tmp_175_fu_1277_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_65_fu_1315_p2 = ((trunc_ln133_31_fu_1287_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_66_fu_1500_p2 = ((tmp_182_fu_1469_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_67_fu_1506_p2 = ((trunc_ln133_32_fu_1479_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_68_fu_1518_p2 = ((tmp_183_fu_1486_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_69_fu_1524_p2 = ((trunc_ln133_33_fu_1496_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_70_fu_1787_p2 = ((tmp_192_fu_1756_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_71_fu_1793_p2 = ((trunc_ln133_34_fu_1766_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_72_fu_1805_p2 = ((tmp_193_fu_1773_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_73_fu_1811_p2 = ((trunc_ln133_35_fu_1783_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_74_fu_2073_p2 = ((tmp_202_fu_2042_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_75_fu_2079_p2 = ((trunc_ln133_36_fu_2052_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_76_fu_2091_p2 = ((tmp_203_fu_2059_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_77_fu_2097_p2 = ((trunc_ln133_37_fu_2069_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_78_fu_2358_p2 = ((tmp_212_fu_2327_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_79_fu_2364_p2 = ((trunc_ln133_38_fu_2337_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_80_fu_2376_p2 = ((tmp_213_fu_2344_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_81_fu_2382_p2 = ((trunc_ln133_39_fu_2354_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_82_fu_2645_p2 = ((tmp_222_fu_2614_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_83_fu_2651_p2 = ((trunc_ln133_40_fu_2624_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_84_fu_2663_p2 = ((tmp_223_fu_2631_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_85_fu_2669_p2 = ((trunc_ln133_41_fu_2641_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_86_fu_2931_p2 = ((tmp_232_fu_2900_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_87_fu_2937_p2 = ((trunc_ln133_42_fu_2910_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_88_fu_2949_p2 = ((tmp_233_fu_2917_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_89_fu_2955_p2 = ((trunc_ln133_43_fu_2927_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_90_fu_3356_p2 = ((tmp_242_fu_3325_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_91_fu_3362_p2 = ((trunc_ln133_44_fu_3335_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_92_fu_3374_p2 = ((tmp_243_fu_3342_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_93_fu_3380_p2 = ((trunc_ln133_45_fu_3352_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_fu_1291_p2 = ((tmp_s_fu_1259_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_27_fu_1722_p2 = ((trunc_ln134_fu_1712_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_28_fu_2003_p2 = ((tmp_195_fu_1989_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_29_fu_2009_p2 = ((trunc_ln134_13_fu_1999_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_30_fu_2288_p2 = ((tmp_205_fu_2274_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_31_fu_2294_p2 = ((trunc_ln134_14_fu_2284_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_32_fu_2574_p2 = ((tmp_215_fu_2560_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_33_fu_2580_p2 = ((trunc_ln134_15_fu_2570_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_34_fu_2861_p2 = ((tmp_225_fu_2847_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_35_fu_2867_p2 = ((trunc_ln134_16_fu_2857_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_36_fu_3146_p2 = ((tmp_235_fu_3132_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_37_fu_3152_p2 = ((trunc_ln134_17_fu_3142_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_38_fu_3427_p2 = ((tmp_245_fu_3413_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_39_fu_3433_p2 = ((trunc_ln134_18_fu_3423_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_fu_1716_p2 = ((tmp_185_fu_1702_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_63_fu_1375_p2 = ((trunc_ln135_fu_1347_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_64_fu_1387_p2 = ((tmp_179_fu_1355_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_65_fu_1393_p2 = ((trunc_ln135_31_fu_1365_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_66_fu_1590_p2 = ((tmp_187_fu_1559_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_67_fu_1596_p2 = ((trunc_ln135_32_fu_1569_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_68_fu_1608_p2 = ((tmp_188_fu_1576_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_69_fu_1614_p2 = ((trunc_ln135_33_fu_1586_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_70_fu_1877_p2 = ((tmp_197_fu_1846_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_71_fu_1883_p2 = ((trunc_ln135_34_fu_1856_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_72_fu_1895_p2 = ((tmp_198_fu_1863_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_73_fu_1901_p2 = ((trunc_ln135_35_fu_1873_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_74_fu_2162_p2 = ((tmp_207_fu_2131_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_75_fu_2168_p2 = ((trunc_ln135_36_fu_2141_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_76_fu_2180_p2 = ((tmp_208_fu_2148_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_77_fu_2186_p2 = ((trunc_ln135_37_fu_2158_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_78_fu_2448_p2 = ((tmp_217_fu_2417_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_79_fu_2454_p2 = ((trunc_ln135_38_fu_2427_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_80_fu_2466_p2 = ((tmp_218_fu_2434_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_81_fu_2472_p2 = ((trunc_ln135_39_fu_2444_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_82_fu_2735_p2 = ((tmp_227_fu_2704_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_83_fu_2741_p2 = ((trunc_ln135_40_fu_2714_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_84_fu_2753_p2 = ((tmp_228_fu_2721_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_85_fu_2759_p2 = ((trunc_ln135_41_fu_2731_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_86_fu_3020_p2 = ((tmp_237_fu_2989_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_87_fu_3026_p2 = ((trunc_ln135_42_fu_2999_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_88_fu_3038_p2 = ((tmp_238_fu_3006_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_89_fu_3044_p2 = ((trunc_ln135_43_fu_3016_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_90_fu_3215_p2 = ((tmp_247_fu_3184_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_91_fu_3221_p2 = ((trunc_ln135_44_fu_3194_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_92_fu_3233_p2 = ((tmp_248_fu_3201_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_93_fu_3239_p2 = ((trunc_ln135_45_fu_3211_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_fu_1369_p2 = ((tmp_178_fu_1337_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_27_fu_1668_p2 = ((trunc_ln136_fu_1658_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_28_fu_1949_p2 = ((tmp_200_fu_1935_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_29_fu_1955_p2 = ((trunc_ln136_13_fu_1945_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_30_fu_2234_p2 = ((tmp_210_fu_2220_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_31_fu_2240_p2 = ((trunc_ln136_14_fu_2230_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_32_fu_2520_p2 = ((tmp_220_fu_2506_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_33_fu_2526_p2 = ((trunc_ln136_15_fu_2516_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_34_fu_2807_p2 = ((tmp_230_fu_2793_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_35_fu_2813_p2 = ((trunc_ln136_16_fu_2803_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_36_fu_3092_p2 = ((tmp_240_fu_3078_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_37_fu_3098_p2 = ((trunc_ln136_17_fu_3088_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_38_fu_3286_p2 = ((tmp_250_fu_3272_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_39_fu_3292_p2 = ((trunc_ln136_18_fu_3282_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_fu_1662_p2 = ((tmp_190_fu_1648_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_11_fu_3503_p2 = ((trunc_ln139_fu_3476_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_12_fu_3515_p2 = ((tmp_253_fu_3483_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_13_fu_3521_p2 = ((trunc_ln139_5_fu_3493_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_14_fu_3556_p2 = ((tmp_255_fu_3542_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_15_fu_3562_p2 = ((trunc_ln139_6_fu_3552_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_fu_3497_p2 = ((tmp_252_fu_3466_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln140_3_fu_3608_p2 = ((trunc_ln140_fu_3598_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln140_fu_3602_p2 = ((tmp_257_fu_3588_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign max1_26_fu_1548_p3 = ((and_ln133_33_fu_1542_p2[0:0] == 1'b1) ? reg_918 : max1_reg_4582);

    assign max1_27_fu_1835_p3 = ((and_ln133_35_fu_1829_p2[0:0] == 1'b1) ? reg_944 : max1_26_reg_4614);

    assign max1_28_fu_2121_p3 = ((and_ln133_37_fu_2115_p2[0:0] == 1'b1) ? n1_39_reg_4596 : max1_27_reg_4647);

    assign max1_29_fu_2406_p3 = ((and_ln133_39_fu_2400_p2[0:0] == 1'b1) ? reg_878 : max1_28_reg_4680);

    assign max1_30_fu_2693_p3 = ((and_ln133_41_fu_2687_p2[0:0] == 1'b1) ? reg_944 : max1_29_reg_4721);

    assign max1_31_fu_2979_p3 = ((and_ln133_43_fu_2973_p2[0:0] == 1'b1) ? n1_48_reg_4708 : max1_30_reg_4772);

    assign max1_32_fu_3404_p3 = ((and_ln133_45_fu_3398_p2[0:0] == 1'b1) ? n1_51_reg_4742 : max1_31_reg_4805);

    assign max1_fu_1443_p3 = ((and_ln133_31_fu_1439_p2[0:0] == 1'b1) ? reg_898 : reg_924);

    assign max2_26_fu_1638_p3 = ((and_ln135_33_fu_1632_p2[0:0] == 1'b1) ? reg_911 : max2_reg_4568);

    assign max2_27_fu_1925_p3 = ((and_ln135_35_fu_1919_p2[0:0] == 1'b1) ? reg_938 : max2_26_reg_4621);

    assign max2_28_fu_2210_p3 = ((and_ln135_37_fu_2204_p2[0:0] == 1'b1) ? reg_930 : max2_27_reg_4654);

    assign max2_29_fu_2496_p3 = ((and_ln135_39_fu_2490_p2[0:0] == 1'b1) ? reg_884 : max2_28_reg_4687);

    assign max2_30_fu_2783_p3 = ((and_ln135_41_fu_2777_p2[0:0] == 1'b1) ? reg_891 : max2_29_reg_4728);

    assign max2_31_fu_3068_p3 = ((and_ln135_43_fu_3062_p2[0:0] == 1'b1) ? reg_938 : max2_30_reg_4779);

    assign max2_32_fu_3263_p3 = ((and_ln135_45_fu_3257_p2[0:0] == 1'b1) ? n2_51_reg_4751 : max2_31_reg_4812);

    assign max2_fu_1417_p3 = ((and_ln135_31_fu_1411_p2[0:0] == 1'b1) ? reg_904 : reg_930);

    assign min1_20_fu_1457_p3 = ((and_ln134_fu_1452_p2[0:0] == 1'b1) ? reg_898 : reg_924);

    assign min1_21_fu_1745_p3 = ((and_ln134_30_fu_1739_p2[0:0] == 1'b1) ? reg_918 : min1_20_reg_4589);

    assign min1_22_fu_2032_p3 = ((and_ln134_32_fu_2026_p2[0:0] == 1'b1) ? reg_944 : min1_21_reg_4635);

    assign min1_23_fu_2317_p3 = ((and_ln134_34_fu_2311_p2[0:0] == 1'b1) ? n1_39_reg_4596 : min1_22_reg_4668);

    assign min1_24_fu_2603_p3 = ((and_ln134_36_fu_2597_p2[0:0] == 1'b1) ? reg_878 : min1_23_reg_4701);

    assign min1_25_fu_2890_p3 = ((and_ln134_38_fu_2884_p2[0:0] == 1'b1) ? reg_944 : min1_24_reg_4760);

    assign min1_26_fu_3175_p3 = ((and_ln134_40_fu_3169_p2[0:0] == 1'b1) ? n1_48_reg_4708 : min1_25_reg_4793);

    assign min1_27_fu_3457_p3 = ((and_ln134_42_fu_3451_p2[0:0] == 1'b1) ? n1_51_reg_4742 : min1_26_reg_4826);

    assign min2_20_fu_1431_p3 = ((and_ln136_fu_1425_p2[0:0] == 1'b1) ? reg_904 : reg_930);

    assign min2_21_fu_1692_p3 = ((and_ln136_30_fu_1686_p2[0:0] == 1'b1) ? reg_911 : min2_20_reg_4575);

    assign min2_22_fu_1979_p3 = ((and_ln136_32_fu_1973_p2[0:0] == 1'b1) ? reg_938 : min2_21_reg_4628);

    assign min2_23_fu_2264_p3 = ((and_ln136_34_fu_2258_p2[0:0] == 1'b1) ? reg_930 : min2_22_reg_4661);

    assign min2_24_fu_2550_p3 = ((and_ln136_36_fu_2544_p2[0:0] == 1'b1) ? reg_884 : min2_23_reg_4694);

    assign min2_25_fu_2837_p3 = ((and_ln136_38_fu_2831_p2[0:0] == 1'b1) ? reg_891 : min2_24_reg_4735);

    assign min2_26_fu_3122_p3 = ((and_ln136_40_fu_3116_p2[0:0] == 1'b1) ? reg_938 : min2_25_reg_4786);

    assign min2_27_fu_3316_p3 = ((and_ln136_42_fu_3310_p2[0:0] == 1'b1) ? n2_51_reg_4751 : min2_26_reg_4819);

    assign mul_ln120_fu_984_p0 = mul_ln120_fu_984_p00;

    assign mul_ln120_fu_984_p00 = p1_offset;

    assign mul_ln120_fu_984_p1 = 7'd27;

    assign or_ln133_31_fu_1321_p2 = (icmp_ln133_65_fu_1315_p2 | icmp_ln133_64_fu_1309_p2);

    assign or_ln133_32_fu_1512_p2 = (icmp_ln133_67_fu_1506_p2 | icmp_ln133_66_fu_1500_p2);

    assign or_ln133_33_fu_1530_p2 = (icmp_ln133_69_fu_1524_p2 | icmp_ln133_68_fu_1518_p2);

    assign or_ln133_34_fu_1799_p2 = (icmp_ln133_71_fu_1793_p2 | icmp_ln133_70_fu_1787_p2);

    assign or_ln133_35_fu_1817_p2 = (icmp_ln133_73_fu_1811_p2 | icmp_ln133_72_fu_1805_p2);

    assign or_ln133_36_fu_2085_p2 = (icmp_ln133_75_fu_2079_p2 | icmp_ln133_74_fu_2073_p2);

    assign or_ln133_37_fu_2103_p2 = (icmp_ln133_77_fu_2097_p2 | icmp_ln133_76_fu_2091_p2);

    assign or_ln133_38_fu_2370_p2 = (icmp_ln133_79_fu_2364_p2 | icmp_ln133_78_fu_2358_p2);

    assign or_ln133_39_fu_2388_p2 = (icmp_ln133_81_fu_2382_p2 | icmp_ln133_80_fu_2376_p2);

    assign or_ln133_40_fu_2657_p2 = (icmp_ln133_83_fu_2651_p2 | icmp_ln133_82_fu_2645_p2);

    assign or_ln133_41_fu_2675_p2 = (icmp_ln133_85_fu_2669_p2 | icmp_ln133_84_fu_2663_p2);

    assign or_ln133_42_fu_2943_p2 = (icmp_ln133_87_fu_2937_p2 | icmp_ln133_86_fu_2931_p2);

    assign or_ln133_43_fu_2961_p2 = (icmp_ln133_89_fu_2955_p2 | icmp_ln133_88_fu_2949_p2);

    assign or_ln133_44_fu_3368_p2 = (icmp_ln133_91_fu_3362_p2 | icmp_ln133_90_fu_3356_p2);

    assign or_ln133_45_fu_3386_p2 = (icmp_ln133_93_fu_3380_p2 | icmp_ln133_92_fu_3374_p2);

    assign or_ln133_fu_1303_p2 = (icmp_ln133_fu_1291_p2 | icmp_ln133_63_fu_1297_p2);

    assign or_ln134_13_fu_2015_p2 = (icmp_ln134_29_fu_2009_p2 | icmp_ln134_28_fu_2003_p2);

    assign or_ln134_14_fu_2300_p2 = (icmp_ln134_31_fu_2294_p2 | icmp_ln134_30_fu_2288_p2);

    assign or_ln134_15_fu_2586_p2 = (icmp_ln134_33_fu_2580_p2 | icmp_ln134_32_fu_2574_p2);

    assign or_ln134_16_fu_2873_p2 = (icmp_ln134_35_fu_2867_p2 | icmp_ln134_34_fu_2861_p2);

    assign or_ln134_17_fu_3158_p2 = (icmp_ln134_37_fu_3152_p2 | icmp_ln134_36_fu_3146_p2);

    assign or_ln134_18_fu_3439_p2 = (icmp_ln134_39_fu_3433_p2 | icmp_ln134_38_fu_3427_p2);

    assign or_ln134_fu_1728_p2 = (icmp_ln134_fu_1716_p2 | icmp_ln134_27_fu_1722_p2);

    assign or_ln135_31_fu_1399_p2 = (icmp_ln135_65_fu_1393_p2 | icmp_ln135_64_fu_1387_p2);

    assign or_ln135_32_fu_1602_p2 = (icmp_ln135_67_fu_1596_p2 | icmp_ln135_66_fu_1590_p2);

    assign or_ln135_33_fu_1620_p2 = (icmp_ln135_69_fu_1614_p2 | icmp_ln135_68_fu_1608_p2);

    assign or_ln135_34_fu_1889_p2 = (icmp_ln135_71_fu_1883_p2 | icmp_ln135_70_fu_1877_p2);

    assign or_ln135_35_fu_1907_p2 = (icmp_ln135_73_fu_1901_p2 | icmp_ln135_72_fu_1895_p2);

    assign or_ln135_36_fu_2174_p2 = (icmp_ln135_75_fu_2168_p2 | icmp_ln135_74_fu_2162_p2);

    assign or_ln135_37_fu_2192_p2 = (icmp_ln135_77_fu_2186_p2 | icmp_ln135_76_fu_2180_p2);

    assign or_ln135_38_fu_2460_p2 = (icmp_ln135_79_fu_2454_p2 | icmp_ln135_78_fu_2448_p2);

    assign or_ln135_39_fu_2478_p2 = (icmp_ln135_81_fu_2472_p2 | icmp_ln135_80_fu_2466_p2);

    assign or_ln135_40_fu_2747_p2 = (icmp_ln135_83_fu_2741_p2 | icmp_ln135_82_fu_2735_p2);

    assign or_ln135_41_fu_2765_p2 = (icmp_ln135_85_fu_2759_p2 | icmp_ln135_84_fu_2753_p2);

    assign or_ln135_42_fu_3032_p2 = (icmp_ln135_87_fu_3026_p2 | icmp_ln135_86_fu_3020_p2);

    assign or_ln135_43_fu_3050_p2 = (icmp_ln135_89_fu_3044_p2 | icmp_ln135_88_fu_3038_p2);

    assign or_ln135_44_fu_3227_p2 = (icmp_ln135_91_fu_3221_p2 | icmp_ln135_90_fu_3215_p2);

    assign or_ln135_45_fu_3245_p2 = (icmp_ln135_93_fu_3239_p2 | icmp_ln135_92_fu_3233_p2);

    assign or_ln135_fu_1381_p2 = (icmp_ln135_fu_1369_p2 | icmp_ln135_63_fu_1375_p2);

    assign or_ln136_13_fu_1961_p2 = (icmp_ln136_29_fu_1955_p2 | icmp_ln136_28_fu_1949_p2);

    assign or_ln136_14_fu_2246_p2 = (icmp_ln136_31_fu_2240_p2 | icmp_ln136_30_fu_2234_p2);

    assign or_ln136_15_fu_2532_p2 = (icmp_ln136_33_fu_2526_p2 | icmp_ln136_32_fu_2520_p2);

    assign or_ln136_16_fu_2819_p2 = (icmp_ln136_35_fu_2813_p2 | icmp_ln136_34_fu_2807_p2);

    assign or_ln136_17_fu_3104_p2 = (icmp_ln136_37_fu_3098_p2 | icmp_ln136_36_fu_3092_p2);

    assign or_ln136_18_fu_3298_p2 = (icmp_ln136_39_fu_3292_p2 | icmp_ln136_38_fu_3286_p2);

    assign or_ln136_fu_1674_p2 = (icmp_ln136_fu_1662_p2 | icmp_ln136_27_fu_1668_p2);

    assign or_ln139_5_fu_3527_p2 = (icmp_ln139_13_fu_3521_p2 | icmp_ln139_12_fu_3515_p2);

    assign or_ln139_6_fu_3568_p2 = (icmp_ln139_15_fu_3562_p2 | icmp_ln139_14_fu_3556_p2);

    assign or_ln139_fu_3509_p2 = (icmp_ln139_fu_3497_p2 | icmp_ln139_11_fu_3503_p2);

    assign or_ln140_7_fu_3614_p2 = (icmp_ln140_fu_3602_p2 | icmp_ln140_3_fu_3608_p2);

    assign or_ln140_8_fu_3669_p2 = (and_ln142_fu_3664_p2 | and_ln140_reg_4899);

    assign or_ln140_fu_3647_p2 = (and_ln141_fu_3642_p2 | and_ln140_12_fu_3637_p2);

    assign p2_0_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_0_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_0_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_1_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_1_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_1_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_2_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_2_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_2_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_3_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_3_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_3_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_4_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_4_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_4_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_5_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_5_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_5_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_6_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_6_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_6_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_7_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_7_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_7_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_8_0_address0 = p2_offset_cast_fu_949_p1;

    assign p2_8_1_address0 = p2_offset_cast_fu_949_p1;

    assign p2_8_2_address0 = p2_offset_cast_fu_949_p1;

    assign p2_offset_cast_fu_949_p1 = p2_offset;

    assign tmp_175_fu_1277_p4 = {{bitcast_ln133_31_fu_1273_p1[62:52]}};

    assign tmp_178_fu_1337_p4 = {{bitcast_ln135_fu_1333_p1[62:52]}};

    assign tmp_179_fu_1355_p4 = {{bitcast_ln135_31_fu_1351_p1[62:52]}};

    assign tmp_182_fu_1469_p4 = {{bitcast_ln133_32_fu_1465_p1[62:52]}};

    assign tmp_183_fu_1486_p4 = {{bitcast_ln133_33_fu_1483_p1[62:52]}};

    assign tmp_185_fu_1702_p4 = {{bitcast_ln134_fu_1699_p1[62:52]}};

    assign tmp_187_fu_1559_p4 = {{bitcast_ln135_32_fu_1555_p1[62:52]}};

    assign tmp_188_fu_1576_p4 = {{bitcast_ln135_33_fu_1573_p1[62:52]}};

    assign tmp_190_fu_1648_p4 = {{bitcast_ln136_fu_1645_p1[62:52]}};

    assign tmp_192_fu_1756_p4 = {{bitcast_ln133_34_fu_1752_p1[62:52]}};

    assign tmp_193_fu_1773_p4 = {{bitcast_ln133_35_fu_1770_p1[62:52]}};

    assign tmp_195_fu_1989_p4 = {{bitcast_ln134_13_fu_1986_p1[62:52]}};

    assign tmp_197_fu_1846_p4 = {{bitcast_ln135_34_fu_1842_p1[62:52]}};

    assign tmp_198_fu_1863_p4 = {{bitcast_ln135_35_fu_1860_p1[62:52]}};

    assign tmp_200_fu_1935_p4 = {{bitcast_ln136_13_fu_1932_p1[62:52]}};

    assign tmp_202_fu_2042_p4 = {{bitcast_ln133_36_fu_2039_p1[62:52]}};

    assign tmp_203_fu_2059_p4 = {{bitcast_ln133_37_fu_2056_p1[62:52]}};

    assign tmp_205_fu_2274_p4 = {{bitcast_ln134_14_fu_2271_p1[62:52]}};

    assign tmp_207_fu_2131_p4 = {{bitcast_ln135_36_fu_2127_p1[62:52]}};

    assign tmp_208_fu_2148_p4 = {{bitcast_ln135_37_fu_2145_p1[62:52]}};

    assign tmp_210_fu_2220_p4 = {{bitcast_ln136_14_fu_2217_p1[62:52]}};

    assign tmp_212_fu_2327_p4 = {{bitcast_ln133_38_fu_2323_p1[62:52]}};

    assign tmp_213_fu_2344_p4 = {{bitcast_ln133_39_fu_2341_p1[62:52]}};

    assign tmp_215_fu_2560_p4 = {{bitcast_ln134_15_fu_2557_p1[62:52]}};

    assign tmp_217_fu_2417_p4 = {{bitcast_ln135_38_fu_2413_p1[62:52]}};

    assign tmp_218_fu_2434_p4 = {{bitcast_ln135_39_fu_2431_p1[62:52]}};

    assign tmp_220_fu_2506_p4 = {{bitcast_ln136_15_fu_2503_p1[62:52]}};

    assign tmp_222_fu_2614_p4 = {{bitcast_ln133_40_fu_2610_p1[62:52]}};

    assign tmp_223_fu_2631_p4 = {{bitcast_ln133_41_fu_2628_p1[62:52]}};

    assign tmp_225_fu_2847_p4 = {{bitcast_ln134_16_fu_2844_p1[62:52]}};

    assign tmp_227_fu_2704_p4 = {{bitcast_ln135_40_fu_2700_p1[62:52]}};

    assign tmp_228_fu_2721_p4 = {{bitcast_ln135_41_fu_2718_p1[62:52]}};

    assign tmp_230_fu_2793_p4 = {{bitcast_ln136_16_fu_2790_p1[62:52]}};

    assign tmp_232_fu_2900_p4 = {{bitcast_ln133_42_fu_2897_p1[62:52]}};

    assign tmp_233_fu_2917_p4 = {{bitcast_ln133_43_fu_2914_p1[62:52]}};

    assign tmp_235_fu_3132_p4 = {{bitcast_ln134_17_fu_3129_p1[62:52]}};

    assign tmp_237_fu_2989_p4 = {{bitcast_ln135_42_fu_2985_p1[62:52]}};

    assign tmp_238_fu_3006_p4 = {{bitcast_ln135_43_fu_3003_p1[62:52]}};

    assign tmp_240_fu_3078_p4 = {{bitcast_ln136_17_fu_3075_p1[62:52]}};

    assign tmp_242_fu_3325_p4 = {{bitcast_ln133_44_fu_3322_p1[62:52]}};

    assign tmp_243_fu_3342_p4 = {{bitcast_ln133_45_fu_3339_p1[62:52]}};

    assign tmp_245_fu_3413_p4 = {{bitcast_ln134_18_fu_3410_p1[62:52]}};

    assign tmp_247_fu_3184_p4 = {{bitcast_ln135_44_fu_3181_p1[62:52]}};

    assign tmp_248_fu_3201_p4 = {{bitcast_ln135_45_fu_3198_p1[62:52]}};

    assign tmp_250_fu_3272_p4 = {{bitcast_ln136_18_fu_3269_p1[62:52]}};

    assign tmp_252_fu_3466_p4 = {{bitcast_ln139_fu_3463_p1[62:52]}};

    assign tmp_253_fu_3483_p4 = {{bitcast_ln139_5_fu_3480_p1[62:52]}};

    assign tmp_255_fu_3542_p4 = {{bitcast_ln139_6_fu_3539_p1[62:52]}};

    assign tmp_257_fu_3588_p4 = {{bitcast_ln140_fu_3585_p1[62:52]}};

    assign tmp_s_fu_1259_p4 = {{bitcast_ln133_fu_1255_p1[62:52]}};

    assign trunc_ln133_31_fu_1287_p1 = bitcast_ln133_31_fu_1273_p1[51:0];

    assign trunc_ln133_32_fu_1479_p1 = bitcast_ln133_32_fu_1465_p1[51:0];

    assign trunc_ln133_33_fu_1496_p1 = bitcast_ln133_33_fu_1483_p1[51:0];

    assign trunc_ln133_34_fu_1766_p1 = bitcast_ln133_34_fu_1752_p1[51:0];

    assign trunc_ln133_35_fu_1783_p1 = bitcast_ln133_35_fu_1770_p1[51:0];

    assign trunc_ln133_36_fu_2052_p1 = bitcast_ln133_36_fu_2039_p1[51:0];

    assign trunc_ln133_37_fu_2069_p1 = bitcast_ln133_37_fu_2056_p1[51:0];

    assign trunc_ln133_38_fu_2337_p1 = bitcast_ln133_38_fu_2323_p1[51:0];

    assign trunc_ln133_39_fu_2354_p1 = bitcast_ln133_39_fu_2341_p1[51:0];

    assign trunc_ln133_40_fu_2624_p1 = bitcast_ln133_40_fu_2610_p1[51:0];

    assign trunc_ln133_41_fu_2641_p1 = bitcast_ln133_41_fu_2628_p1[51:0];

    assign trunc_ln133_42_fu_2910_p1 = bitcast_ln133_42_fu_2897_p1[51:0];

    assign trunc_ln133_43_fu_2927_p1 = bitcast_ln133_43_fu_2914_p1[51:0];

    assign trunc_ln133_44_fu_3335_p1 = bitcast_ln133_44_fu_3322_p1[51:0];

    assign trunc_ln133_45_fu_3352_p1 = bitcast_ln133_45_fu_3339_p1[51:0];

    assign trunc_ln133_fu_1269_p1 = bitcast_ln133_fu_1255_p1[51:0];

    assign trunc_ln134_13_fu_1999_p1 = bitcast_ln134_13_fu_1986_p1[51:0];

    assign trunc_ln134_14_fu_2284_p1 = bitcast_ln134_14_fu_2271_p1[51:0];

    assign trunc_ln134_15_fu_2570_p1 = bitcast_ln134_15_fu_2557_p1[51:0];

    assign trunc_ln134_16_fu_2857_p1 = bitcast_ln134_16_fu_2844_p1[51:0];

    assign trunc_ln134_17_fu_3142_p1 = bitcast_ln134_17_fu_3129_p1[51:0];

    assign trunc_ln134_18_fu_3423_p1 = bitcast_ln134_18_fu_3410_p1[51:0];

    assign trunc_ln134_fu_1712_p1 = bitcast_ln134_fu_1699_p1[51:0];

    assign trunc_ln135_31_fu_1365_p1 = bitcast_ln135_31_fu_1351_p1[51:0];

    assign trunc_ln135_32_fu_1569_p1 = bitcast_ln135_32_fu_1555_p1[51:0];

    assign trunc_ln135_33_fu_1586_p1 = bitcast_ln135_33_fu_1573_p1[51:0];

    assign trunc_ln135_34_fu_1856_p1 = bitcast_ln135_34_fu_1842_p1[51:0];

    assign trunc_ln135_35_fu_1873_p1 = bitcast_ln135_35_fu_1860_p1[51:0];

    assign trunc_ln135_36_fu_2141_p1 = bitcast_ln135_36_fu_2127_p1[51:0];

    assign trunc_ln135_37_fu_2158_p1 = bitcast_ln135_37_fu_2145_p1[51:0];

    assign trunc_ln135_38_fu_2427_p1 = bitcast_ln135_38_fu_2413_p1[51:0];

    assign trunc_ln135_39_fu_2444_p1 = bitcast_ln135_39_fu_2431_p1[51:0];

    assign trunc_ln135_40_fu_2714_p1 = bitcast_ln135_40_fu_2700_p1[51:0];

    assign trunc_ln135_41_fu_2731_p1 = bitcast_ln135_41_fu_2718_p1[51:0];

    assign trunc_ln135_42_fu_2999_p1 = bitcast_ln135_42_fu_2985_p1[51:0];

    assign trunc_ln135_43_fu_3016_p1 = bitcast_ln135_43_fu_3003_p1[51:0];

    assign trunc_ln135_44_fu_3194_p1 = bitcast_ln135_44_fu_3181_p1[51:0];

    assign trunc_ln135_45_fu_3211_p1 = bitcast_ln135_45_fu_3198_p1[51:0];

    assign trunc_ln135_fu_1347_p1 = bitcast_ln135_fu_1333_p1[51:0];

    assign trunc_ln136_13_fu_1945_p1 = bitcast_ln136_13_fu_1932_p1[51:0];

    assign trunc_ln136_14_fu_2230_p1 = bitcast_ln136_14_fu_2217_p1[51:0];

    assign trunc_ln136_15_fu_2516_p1 = bitcast_ln136_15_fu_2503_p1[51:0];

    assign trunc_ln136_16_fu_2803_p1 = bitcast_ln136_16_fu_2790_p1[51:0];

    assign trunc_ln136_17_fu_3088_p1 = bitcast_ln136_17_fu_3075_p1[51:0];

    assign trunc_ln136_18_fu_3282_p1 = bitcast_ln136_18_fu_3269_p1[51:0];

    assign trunc_ln136_fu_1658_p1 = bitcast_ln136_fu_1645_p1[51:0];

    assign trunc_ln139_5_fu_3493_p1 = bitcast_ln139_5_fu_3480_p1[51:0];

    assign trunc_ln139_6_fu_3552_p1 = bitcast_ln139_6_fu_3539_p1[51:0];

    assign trunc_ln139_fu_3476_p1 = bitcast_ln139_fu_3463_p1[51:0];

    assign trunc_ln140_fu_3598_p1 = bitcast_ln140_fu_3585_p1[51:0];

    assign zext_ln120_17_fu_990_p1 = mul_ln120_fu_984_p2;

    assign zext_ln120_18_fu_1040_p1 = add_ln120_fu_1035_p2;

    assign zext_ln120_19_fu_1120_p1 = add_ln120_9_fu_1115_p2;

    assign zext_ln129_47_fu_1050_p1 = add_ln129_47_fu_1045_p2;

    assign zext_ln129_48_fu_1130_p1 = add_ln129_48_fu_1125_p2;

    assign zext_ln129_49_fu_1010_p1 = add_ln129_49_fu_1005_p2;

    assign zext_ln129_50_fu_1060_p1 = add_ln129_50_fu_1055_p2;

    assign zext_ln129_51_fu_1160_p1 = add_ln129_51_fu_1155_p2;

    assign zext_ln129_52_fu_1020_p1 = add_ln129_52_fu_1015_p2;

    assign zext_ln129_53_fu_1080_p1 = add_ln129_53_fu_1075_p2;

    assign zext_ln129_54_fu_1180_p1 = add_ln129_54_fu_1175_p2;

    assign zext_ln129_55_fu_1030_p1 = add_ln129_55_fu_1025_p2;

    assign zext_ln129_56_fu_1100_p1 = add_ln129_56_fu_1095_p2;

    assign zext_ln129_57_fu_1200_p1 = add_ln129_57_fu_1195_p2;

    assign zext_ln129_58_fu_1070_p1 = add_ln129_58_fu_1065_p2;

    assign zext_ln129_59_fu_1140_p1 = add_ln129_59_fu_1135_p2;

    assign zext_ln129_60_fu_1220_p1 = add_ln129_60_fu_1215_p2;

    assign zext_ln129_61_fu_1090_p1 = add_ln129_61_fu_1085_p2;

    assign zext_ln129_62_fu_1170_p1 = add_ln129_62_fu_1165_p2;

    assign zext_ln129_63_fu_1230_p1 = add_ln129_63_fu_1225_p2;

    assign zext_ln129_64_fu_1110_p1 = add_ln129_64_fu_1105_p2;

    assign zext_ln129_65_fu_1190_p1 = add_ln129_65_fu_1185_p2;

    assign zext_ln129_66_fu_1240_p1 = add_ln129_66_fu_1235_p2;

    assign zext_ln129_67_fu_1150_p1 = add_ln129_67_fu_1145_p2;

    assign zext_ln129_68_fu_1210_p1 = add_ln129_68_fu_1205_p2;

    assign zext_ln129_69_fu_1250_p1 = add_ln129_69_fu_1245_p2;

    assign zext_ln129_fu_1000_p1 = add_ln129_fu_995_p2;

endmodule  //main_pointsOverlap_double_s
