/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_forwardKin_Pipeline_VITIS_LOOP_218_3 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    this_TLink_0_0_load,
    this_TLink_0_1_load,
    this_TLink_0_2_load,
    this_TLink_0_3_load,
    this_TLink_1_0_load,
    this_TLink_1_1_load,
    this_TLink_1_2_load,
    this_TLink_1_3_load,
    this_TLink_2_0_load,
    this_TLink_2_1_load,
    this_TLink_2_2_load,
    this_TLink_2_3_load,
    this_TLink_3_0_load,
    this_TLink_3_1_load,
    this_TLink_3_2_load,
    this_TLink_3_3_load,
    this_TJoint_0_0_address0,
    this_TJoint_0_0_ce0,
    this_TJoint_0_0_we0,
    this_TJoint_0_0_d0,
    this_TJoint_0_0_q0,
    this_TJoint_1_0_address0,
    this_TJoint_1_0_ce0,
    this_TJoint_1_0_we0,
    this_TJoint_1_0_d0,
    this_TJoint_1_0_q0,
    this_TJoint_2_0_address0,
    this_TJoint_2_0_ce0,
    this_TJoint_2_0_we0,
    this_TJoint_2_0_d0,
    this_TJoint_2_0_q0,
    this_TJoint_3_0_address0,
    this_TJoint_3_0_ce0,
    this_TJoint_3_0_we0,
    this_TJoint_3_0_d0,
    this_TJoint_3_0_q0,
    this_TCurr_0_0_address0,
    this_TCurr_0_0_ce0,
    this_TCurr_0_0_we0,
    this_TCurr_0_0_d0,
    this_TCurr_0_0_q0,
    this_TJoint_0_1_address0,
    this_TJoint_0_1_ce0,
    this_TJoint_0_1_we0,
    this_TJoint_0_1_d0,
    this_TJoint_0_1_q0,
    this_TJoint_1_1_address0,
    this_TJoint_1_1_ce0,
    this_TJoint_1_1_we0,
    this_TJoint_1_1_d0,
    this_TJoint_1_1_q0,
    this_TJoint_2_1_address0,
    this_TJoint_2_1_ce0,
    this_TJoint_2_1_we0,
    this_TJoint_2_1_d0,
    this_TJoint_2_1_q0,
    this_TJoint_3_1_address0,
    this_TJoint_3_1_ce0,
    this_TJoint_3_1_we0,
    this_TJoint_3_1_d0,
    this_TJoint_3_1_q0,
    this_TCurr_0_1_address0,
    this_TCurr_0_1_ce0,
    this_TCurr_0_1_we0,
    this_TCurr_0_1_d0,
    this_TCurr_0_1_q0,
    this_TJoint_0_2_address0,
    this_TJoint_0_2_ce0,
    this_TJoint_0_2_we0,
    this_TJoint_0_2_d0,
    this_TJoint_0_2_q0,
    this_TJoint_1_2_address0,
    this_TJoint_1_2_ce0,
    this_TJoint_1_2_we0,
    this_TJoint_1_2_d0,
    this_TJoint_1_2_q0,
    this_TJoint_2_2_address0,
    this_TJoint_2_2_ce0,
    this_TJoint_2_2_we0,
    this_TJoint_2_2_d0,
    this_TJoint_2_2_q0,
    this_TJoint_3_2_address0,
    this_TJoint_3_2_ce0,
    this_TJoint_3_2_we0,
    this_TJoint_3_2_d0,
    this_TJoint_3_2_q0,
    this_TCurr_0_2_address0,
    this_TCurr_0_2_ce0,
    this_TCurr_0_2_we0,
    this_TCurr_0_2_d0,
    this_TCurr_0_2_q0,
    this_TJoint_0_3_address0,
    this_TJoint_0_3_ce0,
    this_TJoint_0_3_we0,
    this_TJoint_0_3_d0,
    this_TJoint_0_3_q0,
    this_TJoint_1_3_address0,
    this_TJoint_1_3_ce0,
    this_TJoint_1_3_we0,
    this_TJoint_1_3_d0,
    this_TJoint_1_3_q0,
    this_TJoint_2_3_address0,
    this_TJoint_2_3_ce0,
    this_TJoint_2_3_we0,
    this_TJoint_2_3_d0,
    this_TJoint_2_3_q0,
    this_TJoint_3_3_address0,
    this_TJoint_3_3_ce0,
    this_TJoint_3_3_we0,
    this_TJoint_3_3_d0,
    this_TJoint_3_3_q0,
    this_TCurr_0_3_address0,
    this_TCurr_0_3_ce0,
    this_TCurr_0_3_we0,
    this_TCurr_0_3_d0,
    this_TCurr_0_3_q0,
    this_TCurr_1_0_address0,
    this_TCurr_1_0_ce0,
    this_TCurr_1_0_we0,
    this_TCurr_1_0_d0,
    this_TCurr_1_0_q0,
    this_TCurr_1_1_address0,
    this_TCurr_1_1_ce0,
    this_TCurr_1_1_we0,
    this_TCurr_1_1_d0,
    this_TCurr_1_1_q0,
    this_TCurr_1_2_address0,
    this_TCurr_1_2_ce0,
    this_TCurr_1_2_we0,
    this_TCurr_1_2_d0,
    this_TCurr_1_2_q0,
    this_TCurr_1_3_address0,
    this_TCurr_1_3_ce0,
    this_TCurr_1_3_we0,
    this_TCurr_1_3_d0,
    this_TCurr_1_3_q0,
    this_TCurr_2_0_address0,
    this_TCurr_2_0_ce0,
    this_TCurr_2_0_we0,
    this_TCurr_2_0_d0,
    this_TCurr_2_0_q0,
    this_TCurr_2_1_address0,
    this_TCurr_2_1_ce0,
    this_TCurr_2_1_we0,
    this_TCurr_2_1_d0,
    this_TCurr_2_1_q0,
    this_TCurr_2_2_address0,
    this_TCurr_2_2_ce0,
    this_TCurr_2_2_we0,
    this_TCurr_2_2_d0,
    this_TCurr_2_2_q0,
    this_TCurr_2_3_address0,
    this_TCurr_2_3_ce0,
    this_TCurr_2_3_we0,
    this_TCurr_2_3_d0,
    this_TCurr_2_3_q0,
    this_TCurr_3_0_address0,
    this_TCurr_3_0_ce0,
    this_TCurr_3_0_we0,
    this_TCurr_3_0_d0,
    this_TCurr_3_0_q0,
    this_TCurr_3_1_address0,
    this_TCurr_3_1_ce0,
    this_TCurr_3_1_we0,
    this_TCurr_3_1_d0,
    this_TCurr_3_1_q0,
    this_TCurr_3_2_address0,
    this_TCurr_3_2_ce0,
    this_TCurr_3_2_we0,
    this_TCurr_3_2_d0,
    this_TCurr_3_2_q0,
    this_TCurr_3_3_address0,
    this_TCurr_3_3_ce0,
    this_TCurr_3_3_we0,
    this_TCurr_3_3_d0,
    this_TCurr_3_3_q0,
    this_q_address0,
    this_q_ce0,
    this_q_q0,
    this_TLink_0_0_address0,
    this_TLink_0_0_ce0,
    this_TLink_0_0_q0,
    this_TLink_1_0_address0,
    this_TLink_1_0_ce0,
    this_TLink_1_0_q0,
    this_TLink_2_0_address0,
    this_TLink_2_0_ce0,
    this_TLink_2_0_q0,
    this_TLink_3_0_address0,
    this_TLink_3_0_ce0,
    this_TLink_3_0_q0,
    this_TLink_0_1_address0,
    this_TLink_0_1_ce0,
    this_TLink_0_1_q0,
    this_TLink_1_1_address0,
    this_TLink_1_1_ce0,
    this_TLink_1_1_q0,
    this_TLink_2_1_address0,
    this_TLink_2_1_ce0,
    this_TLink_2_1_q0,
    this_TLink_3_1_address0,
    this_TLink_3_1_ce0,
    this_TLink_3_1_q0,
    this_TLink_0_2_address0,
    this_TLink_0_2_ce0,
    this_TLink_0_2_q0,
    this_TLink_1_2_address0,
    this_TLink_1_2_ce0,
    this_TLink_1_2_q0,
    this_TLink_2_2_address0,
    this_TLink_2_2_ce0,
    this_TLink_2_2_q0,
    this_TLink_3_2_address0,
    this_TLink_3_2_ce0,
    this_TLink_3_2_q0,
    this_TLink_0_3_address0,
    this_TLink_0_3_ce0,
    this_TLink_0_3_q0,
    this_TLink_1_3_address0,
    this_TLink_1_3_ce0,
    this_TLink_1_3_q0,
    this_TLink_2_3_address0,
    this_TLink_2_3_ce0,
    this_TLink_2_3_q0,
    this_TLink_3_3_address0,
    this_TLink_3_3_ce0,
    this_TLink_3_3_q0
);

    parameter ap_ST_fsm_pp0_stage0 = 73'd1;
    parameter ap_ST_fsm_pp0_stage1 = 73'd2;
    parameter ap_ST_fsm_pp0_stage2 = 73'd4;
    parameter ap_ST_fsm_pp0_stage3 = 73'd8;
    parameter ap_ST_fsm_pp0_stage4 = 73'd16;
    parameter ap_ST_fsm_pp0_stage5 = 73'd32;
    parameter ap_ST_fsm_pp0_stage6 = 73'd64;
    parameter ap_ST_fsm_pp0_stage7 = 73'd128;
    parameter ap_ST_fsm_pp0_stage8 = 73'd256;
    parameter ap_ST_fsm_pp0_stage9 = 73'd512;
    parameter ap_ST_fsm_pp0_stage10 = 73'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 73'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 73'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 73'd8192;
    parameter ap_ST_fsm_pp0_stage14 = 73'd16384;
    parameter ap_ST_fsm_pp0_stage15 = 73'd32768;
    parameter ap_ST_fsm_pp0_stage16 = 73'd65536;
    parameter ap_ST_fsm_pp0_stage17 = 73'd131072;
    parameter ap_ST_fsm_pp0_stage18 = 73'd262144;
    parameter ap_ST_fsm_pp0_stage19 = 73'd524288;
    parameter ap_ST_fsm_pp0_stage20 = 73'd1048576;
    parameter ap_ST_fsm_pp0_stage21 = 73'd2097152;
    parameter ap_ST_fsm_pp0_stage22 = 73'd4194304;
    parameter ap_ST_fsm_pp0_stage23 = 73'd8388608;
    parameter ap_ST_fsm_pp0_stage24 = 73'd16777216;
    parameter ap_ST_fsm_pp0_stage25 = 73'd33554432;
    parameter ap_ST_fsm_pp0_stage26 = 73'd67108864;
    parameter ap_ST_fsm_pp0_stage27 = 73'd134217728;
    parameter ap_ST_fsm_pp0_stage28 = 73'd268435456;
    parameter ap_ST_fsm_pp0_stage29 = 73'd536870912;
    parameter ap_ST_fsm_pp0_stage30 = 73'd1073741824;
    parameter ap_ST_fsm_pp0_stage31 = 73'd2147483648;
    parameter ap_ST_fsm_pp0_stage32 = 73'd4294967296;
    parameter ap_ST_fsm_pp0_stage33 = 73'd8589934592;
    parameter ap_ST_fsm_pp0_stage34 = 73'd17179869184;
    parameter ap_ST_fsm_pp0_stage35 = 73'd34359738368;
    parameter ap_ST_fsm_pp0_stage36 = 73'd68719476736;
    parameter ap_ST_fsm_pp0_stage37 = 73'd137438953472;
    parameter ap_ST_fsm_pp0_stage38 = 73'd274877906944;
    parameter ap_ST_fsm_pp0_stage39 = 73'd549755813888;
    parameter ap_ST_fsm_pp0_stage40 = 73'd1099511627776;
    parameter ap_ST_fsm_pp0_stage41 = 73'd2199023255552;
    parameter ap_ST_fsm_pp0_stage42 = 73'd4398046511104;
    parameter ap_ST_fsm_pp0_stage43 = 73'd8796093022208;
    parameter ap_ST_fsm_pp0_stage44 = 73'd17592186044416;
    parameter ap_ST_fsm_pp0_stage45 = 73'd35184372088832;
    parameter ap_ST_fsm_pp0_stage46 = 73'd70368744177664;
    parameter ap_ST_fsm_pp0_stage47 = 73'd140737488355328;
    parameter ap_ST_fsm_pp0_stage48 = 73'd281474976710656;
    parameter ap_ST_fsm_pp0_stage49 = 73'd562949953421312;
    parameter ap_ST_fsm_pp0_stage50 = 73'd1125899906842624;
    parameter ap_ST_fsm_pp0_stage51 = 73'd2251799813685248;
    parameter ap_ST_fsm_pp0_stage52 = 73'd4503599627370496;
    parameter ap_ST_fsm_pp0_stage53 = 73'd9007199254740992;
    parameter ap_ST_fsm_pp0_stage54 = 73'd18014398509481984;
    parameter ap_ST_fsm_pp0_stage55 = 73'd36028797018963968;
    parameter ap_ST_fsm_pp0_stage56 = 73'd72057594037927936;
    parameter ap_ST_fsm_pp0_stage57 = 73'd144115188075855872;
    parameter ap_ST_fsm_pp0_stage58 = 73'd288230376151711744;
    parameter ap_ST_fsm_pp0_stage59 = 73'd576460752303423488;
    parameter ap_ST_fsm_pp0_stage60 = 73'd1152921504606846976;
    parameter ap_ST_fsm_pp0_stage61 = 73'd2305843009213693952;
    parameter ap_ST_fsm_pp0_stage62 = 73'd4611686018427387904;
    parameter ap_ST_fsm_pp0_stage63 = 73'd9223372036854775808;
    parameter ap_ST_fsm_pp0_stage64 = 73'd18446744073709551616;
    parameter ap_ST_fsm_pp0_stage65 = 73'd36893488147419103232;
    parameter ap_ST_fsm_pp0_stage66 = 73'd73786976294838206464;
    parameter ap_ST_fsm_pp0_stage67 = 73'd147573952589676412928;
    parameter ap_ST_fsm_pp0_stage68 = 73'd295147905179352825856;
    parameter ap_ST_fsm_pp0_stage69 = 73'd590295810358705651712;
    parameter ap_ST_fsm_pp0_stage70 = 73'd1180591620717411303424;
    parameter ap_ST_fsm_pp0_stage71 = 73'd2361183241434822606848;
    parameter ap_ST_fsm_pp0_stage72 = 73'd4722366482869645213696;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] this_TLink_0_0_load;
    input [63:0] this_TLink_0_1_load;
    input [63:0] this_TLink_0_2_load;
    input [63:0] this_TLink_0_3_load;
    input [63:0] this_TLink_1_0_load;
    input [63:0] this_TLink_1_1_load;
    input [63:0] this_TLink_1_2_load;
    input [63:0] this_TLink_1_3_load;
    input [63:0] this_TLink_2_0_load;
    input [63:0] this_TLink_2_1_load;
    input [63:0] this_TLink_2_2_load;
    input [63:0] this_TLink_2_3_load;
    input [63:0] this_TLink_3_0_load;
    input [63:0] this_TLink_3_1_load;
    input [63:0] this_TLink_3_2_load;
    input [63:0] this_TLink_3_3_load;
    output [2:0] this_TJoint_0_0_address0;
    output this_TJoint_0_0_ce0;
    output this_TJoint_0_0_we0;
    output [63:0] this_TJoint_0_0_d0;
    input [63:0] this_TJoint_0_0_q0;
    output [2:0] this_TJoint_1_0_address0;
    output this_TJoint_1_0_ce0;
    output this_TJoint_1_0_we0;
    output [63:0] this_TJoint_1_0_d0;
    input [63:0] this_TJoint_1_0_q0;
    output [2:0] this_TJoint_2_0_address0;
    output this_TJoint_2_0_ce0;
    output this_TJoint_2_0_we0;
    output [63:0] this_TJoint_2_0_d0;
    input [63:0] this_TJoint_2_0_q0;
    output [2:0] this_TJoint_3_0_address0;
    output this_TJoint_3_0_ce0;
    output this_TJoint_3_0_we0;
    output [63:0] this_TJoint_3_0_d0;
    input [63:0] this_TJoint_3_0_q0;
    output [2:0] this_TCurr_0_0_address0;
    output this_TCurr_0_0_ce0;
    output this_TCurr_0_0_we0;
    output [63:0] this_TCurr_0_0_d0;
    input [63:0] this_TCurr_0_0_q0;
    output [2:0] this_TJoint_0_1_address0;
    output this_TJoint_0_1_ce0;
    output this_TJoint_0_1_we0;
    output [63:0] this_TJoint_0_1_d0;
    input [63:0] this_TJoint_0_1_q0;
    output [2:0] this_TJoint_1_1_address0;
    output this_TJoint_1_1_ce0;
    output this_TJoint_1_1_we0;
    output [63:0] this_TJoint_1_1_d0;
    input [63:0] this_TJoint_1_1_q0;
    output [2:0] this_TJoint_2_1_address0;
    output this_TJoint_2_1_ce0;
    output this_TJoint_2_1_we0;
    output [63:0] this_TJoint_2_1_d0;
    input [63:0] this_TJoint_2_1_q0;
    output [2:0] this_TJoint_3_1_address0;
    output this_TJoint_3_1_ce0;
    output this_TJoint_3_1_we0;
    output [63:0] this_TJoint_3_1_d0;
    input [63:0] this_TJoint_3_1_q0;
    output [2:0] this_TCurr_0_1_address0;
    output this_TCurr_0_1_ce0;
    output this_TCurr_0_1_we0;
    output [63:0] this_TCurr_0_1_d0;
    input [63:0] this_TCurr_0_1_q0;
    output [2:0] this_TJoint_0_2_address0;
    output this_TJoint_0_2_ce0;
    output this_TJoint_0_2_we0;
    output [63:0] this_TJoint_0_2_d0;
    input [63:0] this_TJoint_0_2_q0;
    output [2:0] this_TJoint_1_2_address0;
    output this_TJoint_1_2_ce0;
    output this_TJoint_1_2_we0;
    output [63:0] this_TJoint_1_2_d0;
    input [63:0] this_TJoint_1_2_q0;
    output [2:0] this_TJoint_2_2_address0;
    output this_TJoint_2_2_ce0;
    output this_TJoint_2_2_we0;
    output [63:0] this_TJoint_2_2_d0;
    input [63:0] this_TJoint_2_2_q0;
    output [2:0] this_TJoint_3_2_address0;
    output this_TJoint_3_2_ce0;
    output this_TJoint_3_2_we0;
    output [63:0] this_TJoint_3_2_d0;
    input [63:0] this_TJoint_3_2_q0;
    output [2:0] this_TCurr_0_2_address0;
    output this_TCurr_0_2_ce0;
    output this_TCurr_0_2_we0;
    output [63:0] this_TCurr_0_2_d0;
    input [63:0] this_TCurr_0_2_q0;
    output [2:0] this_TJoint_0_3_address0;
    output this_TJoint_0_3_ce0;
    output this_TJoint_0_3_we0;
    output [63:0] this_TJoint_0_3_d0;
    input [63:0] this_TJoint_0_3_q0;
    output [2:0] this_TJoint_1_3_address0;
    output this_TJoint_1_3_ce0;
    output this_TJoint_1_3_we0;
    output [63:0] this_TJoint_1_3_d0;
    input [63:0] this_TJoint_1_3_q0;
    output [2:0] this_TJoint_2_3_address0;
    output this_TJoint_2_3_ce0;
    output this_TJoint_2_3_we0;
    output [63:0] this_TJoint_2_3_d0;
    input [63:0] this_TJoint_2_3_q0;
    output [2:0] this_TJoint_3_3_address0;
    output this_TJoint_3_3_ce0;
    output this_TJoint_3_3_we0;
    output [63:0] this_TJoint_3_3_d0;
    input [63:0] this_TJoint_3_3_q0;
    output [2:0] this_TCurr_0_3_address0;
    output this_TCurr_0_3_ce0;
    output this_TCurr_0_3_we0;
    output [63:0] this_TCurr_0_3_d0;
    input [63:0] this_TCurr_0_3_q0;
    output [2:0] this_TCurr_1_0_address0;
    output this_TCurr_1_0_ce0;
    output this_TCurr_1_0_we0;
    output [63:0] this_TCurr_1_0_d0;
    input [63:0] this_TCurr_1_0_q0;
    output [2:0] this_TCurr_1_1_address0;
    output this_TCurr_1_1_ce0;
    output this_TCurr_1_1_we0;
    output [63:0] this_TCurr_1_1_d0;
    input [63:0] this_TCurr_1_1_q0;
    output [2:0] this_TCurr_1_2_address0;
    output this_TCurr_1_2_ce0;
    output this_TCurr_1_2_we0;
    output [63:0] this_TCurr_1_2_d0;
    input [63:0] this_TCurr_1_2_q0;
    output [2:0] this_TCurr_1_3_address0;
    output this_TCurr_1_3_ce0;
    output this_TCurr_1_3_we0;
    output [63:0] this_TCurr_1_3_d0;
    input [63:0] this_TCurr_1_3_q0;
    output [2:0] this_TCurr_2_0_address0;
    output this_TCurr_2_0_ce0;
    output this_TCurr_2_0_we0;
    output [63:0] this_TCurr_2_0_d0;
    input [63:0] this_TCurr_2_0_q0;
    output [2:0] this_TCurr_2_1_address0;
    output this_TCurr_2_1_ce0;
    output this_TCurr_2_1_we0;
    output [63:0] this_TCurr_2_1_d0;
    input [63:0] this_TCurr_2_1_q0;
    output [2:0] this_TCurr_2_2_address0;
    output this_TCurr_2_2_ce0;
    output this_TCurr_2_2_we0;
    output [63:0] this_TCurr_2_2_d0;
    input [63:0] this_TCurr_2_2_q0;
    output [2:0] this_TCurr_2_3_address0;
    output this_TCurr_2_3_ce0;
    output this_TCurr_2_3_we0;
    output [63:0] this_TCurr_2_3_d0;
    input [63:0] this_TCurr_2_3_q0;
    output [2:0] this_TCurr_3_0_address0;
    output this_TCurr_3_0_ce0;
    output this_TCurr_3_0_we0;
    output [63:0] this_TCurr_3_0_d0;
    input [63:0] this_TCurr_3_0_q0;
    output [2:0] this_TCurr_3_1_address0;
    output this_TCurr_3_1_ce0;
    output this_TCurr_3_1_we0;
    output [63:0] this_TCurr_3_1_d0;
    input [63:0] this_TCurr_3_1_q0;
    output [2:0] this_TCurr_3_2_address0;
    output this_TCurr_3_2_ce0;
    output this_TCurr_3_2_we0;
    output [63:0] this_TCurr_3_2_d0;
    input [63:0] this_TCurr_3_2_q0;
    output [2:0] this_TCurr_3_3_address0;
    output this_TCurr_3_3_ce0;
    output this_TCurr_3_3_we0;
    output [63:0] this_TCurr_3_3_d0;
    input [63:0] this_TCurr_3_3_q0;
    output [2:0] this_q_address0;
    output this_q_ce0;
    input [63:0] this_q_q0;
    output [2:0] this_TLink_0_0_address0;
    output this_TLink_0_0_ce0;
    input [63:0] this_TLink_0_0_q0;
    output [2:0] this_TLink_1_0_address0;
    output this_TLink_1_0_ce0;
    input [63:0] this_TLink_1_0_q0;
    output [2:0] this_TLink_2_0_address0;
    output this_TLink_2_0_ce0;
    input [63:0] this_TLink_2_0_q0;
    output [2:0] this_TLink_3_0_address0;
    output this_TLink_3_0_ce0;
    input [63:0] this_TLink_3_0_q0;
    output [2:0] this_TLink_0_1_address0;
    output this_TLink_0_1_ce0;
    input [63:0] this_TLink_0_1_q0;
    output [2:0] this_TLink_1_1_address0;
    output this_TLink_1_1_ce0;
    input [63:0] this_TLink_1_1_q0;
    output [2:0] this_TLink_2_1_address0;
    output this_TLink_2_1_ce0;
    input [63:0] this_TLink_2_1_q0;
    output [2:0] this_TLink_3_1_address0;
    output this_TLink_3_1_ce0;
    input [63:0] this_TLink_3_1_q0;
    output [2:0] this_TLink_0_2_address0;
    output this_TLink_0_2_ce0;
    input [63:0] this_TLink_0_2_q0;
    output [2:0] this_TLink_1_2_address0;
    output this_TLink_1_2_ce0;
    input [63:0] this_TLink_1_2_q0;
    output [2:0] this_TLink_2_2_address0;
    output this_TLink_2_2_ce0;
    input [63:0] this_TLink_2_2_q0;
    output [2:0] this_TLink_3_2_address0;
    output this_TLink_3_2_ce0;
    input [63:0] this_TLink_3_2_q0;
    output [2:0] this_TLink_0_3_address0;
    output this_TLink_0_3_ce0;
    input [63:0] this_TLink_0_3_q0;
    output [2:0] this_TLink_1_3_address0;
    output this_TLink_1_3_ce0;
    input [63:0] this_TLink_1_3_q0;
    output [2:0] this_TLink_2_3_address0;
    output this_TLink_2_3_ce0;
    input [63:0] this_TLink_2_3_q0;
    output [2:0] this_TLink_3_3_address0;
    output this_TLink_3_3_ce0;
    input [63:0] this_TLink_3_3_q0;

    reg ap_idle;
    reg[2:0] this_TJoint_0_0_address0;
    reg this_TJoint_0_0_ce0;
    reg this_TJoint_0_0_we0;
    reg[63:0] this_TJoint_0_0_d0;
    reg[2:0] this_TJoint_1_0_address0;
    reg this_TJoint_1_0_ce0;
    reg this_TJoint_1_0_we0;
    reg[63:0] this_TJoint_1_0_d0;
    reg[2:0] this_TJoint_2_0_address0;
    reg this_TJoint_2_0_ce0;
    reg this_TJoint_2_0_we0;
    reg[63:0] this_TJoint_2_0_d0;
    reg[2:0] this_TJoint_3_0_address0;
    reg this_TJoint_3_0_ce0;
    reg this_TJoint_3_0_we0;
    reg[2:0] this_TCurr_0_0_address0;
    reg this_TCurr_0_0_ce0;
    reg this_TCurr_0_0_we0;
    reg[2:0] this_TJoint_0_1_address0;
    reg this_TJoint_0_1_ce0;
    reg this_TJoint_0_1_we0;
    reg[63:0] this_TJoint_0_1_d0;
    reg[2:0] this_TJoint_1_1_address0;
    reg this_TJoint_1_1_ce0;
    reg this_TJoint_1_1_we0;
    reg[63:0] this_TJoint_1_1_d0;
    reg[2:0] this_TJoint_2_1_address0;
    reg this_TJoint_2_1_ce0;
    reg this_TJoint_2_1_we0;
    reg[63:0] this_TJoint_2_1_d0;
    reg[2:0] this_TJoint_3_1_address0;
    reg this_TJoint_3_1_ce0;
    reg this_TJoint_3_1_we0;
    reg[2:0] this_TCurr_0_1_address0;
    reg this_TCurr_0_1_ce0;
    reg this_TCurr_0_1_we0;
    reg[63:0] this_TCurr_0_1_d0;
    reg[2:0] this_TJoint_0_2_address0;
    reg this_TJoint_0_2_ce0;
    reg this_TJoint_0_2_we0;
    reg[63:0] this_TJoint_0_2_d0;
    reg[2:0] this_TJoint_1_2_address0;
    reg this_TJoint_1_2_ce0;
    reg this_TJoint_1_2_we0;
    reg[63:0] this_TJoint_1_2_d0;
    reg[2:0] this_TJoint_2_2_address0;
    reg this_TJoint_2_2_ce0;
    reg this_TJoint_2_2_we0;
    reg[63:0] this_TJoint_2_2_d0;
    reg[2:0] this_TJoint_3_2_address0;
    reg this_TJoint_3_2_ce0;
    reg this_TJoint_3_2_we0;
    reg[2:0] this_TCurr_0_2_address0;
    reg this_TCurr_0_2_ce0;
    reg this_TCurr_0_2_we0;
    reg[2:0] this_TJoint_0_3_address0;
    reg this_TJoint_0_3_ce0;
    reg this_TJoint_0_3_we0;
    reg[2:0] this_TJoint_1_3_address0;
    reg this_TJoint_1_3_ce0;
    reg this_TJoint_1_3_we0;
    reg[2:0] this_TJoint_2_3_address0;
    reg this_TJoint_2_3_ce0;
    reg this_TJoint_2_3_we0;
    reg[2:0] this_TJoint_3_3_address0;
    reg this_TJoint_3_3_ce0;
    reg this_TJoint_3_3_we0;
    reg[2:0] this_TCurr_0_3_address0;
    reg this_TCurr_0_3_ce0;
    reg this_TCurr_0_3_we0;
    reg[63:0] this_TCurr_0_3_d0;
    reg[2:0] this_TCurr_1_0_address0;
    reg this_TCurr_1_0_ce0;
    reg this_TCurr_1_0_we0;
    reg[63:0] this_TCurr_1_0_d0;
    reg[2:0] this_TCurr_1_1_address0;
    reg this_TCurr_1_1_ce0;
    reg this_TCurr_1_1_we0;
    reg[63:0] this_TCurr_1_1_d0;
    reg[2:0] this_TCurr_1_2_address0;
    reg this_TCurr_1_2_ce0;
    reg this_TCurr_1_2_we0;
    reg[2:0] this_TCurr_1_3_address0;
    reg this_TCurr_1_3_ce0;
    reg this_TCurr_1_3_we0;
    reg[63:0] this_TCurr_1_3_d0;
    reg[2:0] this_TCurr_2_0_address0;
    reg this_TCurr_2_0_ce0;
    reg this_TCurr_2_0_we0;
    reg[63:0] this_TCurr_2_0_d0;
    reg[2:0] this_TCurr_2_1_address0;
    reg this_TCurr_2_1_ce0;
    reg this_TCurr_2_1_we0;
    reg[63:0] this_TCurr_2_1_d0;
    reg[2:0] this_TCurr_2_2_address0;
    reg this_TCurr_2_2_ce0;
    reg this_TCurr_2_2_we0;
    reg[2:0] this_TCurr_2_3_address0;
    reg this_TCurr_2_3_ce0;
    reg this_TCurr_2_3_we0;
    reg[63:0] this_TCurr_2_3_d0;
    reg[2:0] this_TCurr_3_0_address0;
    reg this_TCurr_3_0_ce0;
    reg this_TCurr_3_0_we0;
    reg[63:0] this_TCurr_3_0_d0;
    reg[2:0] this_TCurr_3_1_address0;
    reg this_TCurr_3_1_ce0;
    reg this_TCurr_3_1_we0;
    reg[63:0] this_TCurr_3_1_d0;
    reg[2:0] this_TCurr_3_2_address0;
    reg this_TCurr_3_2_ce0;
    reg this_TCurr_3_2_we0;
    reg[2:0] this_TCurr_3_3_address0;
    reg this_TCurr_3_3_ce0;
    reg this_TCurr_3_3_we0;
    reg[63:0] this_TCurr_3_3_d0;
    reg[2:0] this_q_address0;
    reg this_q_ce0;
    reg this_TLink_0_0_ce0;
    reg this_TLink_1_0_ce0;
    reg this_TLink_2_0_ce0;
    reg this_TLink_3_0_ce0;
    reg this_TLink_0_1_ce0;
    reg this_TLink_1_1_ce0;
    reg this_TLink_2_1_ce0;
    reg this_TLink_3_1_ce0;
    reg this_TLink_0_2_ce0;
    reg this_TLink_1_2_ce0;
    reg this_TLink_2_2_ce0;
    reg this_TLink_3_2_ce0;
    reg this_TLink_0_3_ce0;
    reg this_TLink_1_3_ce0;
    reg this_TLink_2_3_ce0;
    reg this_TLink_3_3_ce0;

    (* fsm_encoding = "none" *) reg   [72:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage23;
    wire    ap_block_pp0_stage23_subdone;
    reg   [0:0] icmp_ln218_reg_3292;
    reg    ap_condition_exit_pp0_iter0_stage23;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_CS_fsm_pp0_stage72;
    wire    ap_block_pp0_stage72_subdone;
    wire   [2:0] l_axis_0_address0;
    reg    l_axis_0_ce0;
    wire   [63:0] l_axis_0_q0;
    reg   [2:0] l_axis_1_address0;
    reg    l_axis_1_ce0;
    wire   [63:0] l_axis_1_q0;
    reg   [2:0] l_axis_2_address0;
    reg    l_axis_2_ce0;
    wire   [63:0] l_axis_2_q0;
    reg   [63:0] reg_1977;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    wire    ap_CS_fsm_pp0_stage17;
    wire    ap_block_pp0_stage17_11001;
    reg   [63:0] reg_1982;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire    ap_CS_fsm_pp0_stage14;
    wire    ap_block_pp0_stage14_11001;
    wire    ap_CS_fsm_pp0_stage20;
    wire    ap_block_pp0_stage20_11001;
    reg   [63:0] reg_1987;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    wire    ap_block_pp0_stage23_11001;
    reg   [63:0] reg_1992;
    wire    ap_CS_fsm_pp0_stage25;
    wire    ap_block_pp0_stage25_11001;
    reg   [0:0] icmp_ln263_reg_3394;
    reg   [63:0] reg_1999;
    reg   [63:0] reg_2006;
    reg   [63:0] reg_2013;
    reg   [63:0] reg_2025;
    reg   [63:0] reg_2035;
    reg   [63:0] reg_2045;
    wire   [63:0] grp_fu_1922_p2;
    reg   [63:0] reg_2052;
    wire    ap_CS_fsm_pp0_stage31;
    wire    ap_block_pp0_stage31_11001;
    wire    ap_CS_fsm_pp0_stage54;
    wire    ap_block_pp0_stage54_11001;
    wire   [63:0] grp_fu_1926_p2;
    reg   [63:0] reg_2058;
    wire    ap_CS_fsm_pp0_stage61;
    wire    ap_block_pp0_stage61_11001;
    wire   [63:0] grp_fu_1930_p2;
    reg   [63:0] reg_2064;
    wire   [63:0] grp_fu_1934_p2;
    reg   [63:0] reg_2070;
    wire   [63:0] grp_fu_1938_p2;
    reg   [63:0] reg_2077;
    wire   [63:0] grp_fu_1942_p2;
    reg   [63:0] reg_2082;
    wire   [63:0] grp_fu_1946_p2;
    reg   [63:0] reg_2089;
    wire   [63:0] grp_fu_1950_p2;
    reg   [63:0] reg_2095;
    wire   [63:0] grp_fu_1954_p2;
    reg   [63:0] reg_2102;
    wire    ap_CS_fsm_pp0_stage66;
    wire    ap_block_pp0_stage66_11001;
    wire   [63:0] grp_fu_1958_p2;
    reg   [63:0] reg_2108;
    wire   [63:0] grp_fu_1962_p2;
    reg   [63:0] reg_2114;
    wire   [63:0] grp_fu_1966_p2;
    reg   [63:0] reg_2120;
    reg   [63:0] reg_2126;
    wire    ap_CS_fsm_pp0_stage32;
    wire    ap_block_pp0_stage32_11001;
    wire    ap_CS_fsm_pp0_stage60;
    wire    ap_block_pp0_stage60_11001;
    wire    ap_CS_fsm_pp0_stage68;
    wire    ap_block_pp0_stage68_11001;
    reg   [63:0] reg_2132;
    reg   [63:0] reg_2138;
    reg   [63:0] reg_2145;
    reg   [63:0] reg_2152;
    reg   [63:0] reg_2159;
    reg   [63:0] reg_2167;
    reg   [63:0] reg_2174;
    reg   [63:0] reg_2182;
    wire    ap_CS_fsm_pp0_stage67;
    wire    ap_block_pp0_stage67_11001;
    reg   [63:0] reg_2189;
    reg   [63:0] reg_2196;
    reg   [63:0] reg_2203;
    reg   [63:0] reg_2209;
    wire    ap_CS_fsm_pp0_stage33;
    wire    ap_block_pp0_stage33_11001;
    reg   [63:0] reg_2214;
    reg   [63:0] reg_2220;
    reg   [63:0] reg_2225;
    reg   [63:0] reg_2233;
    reg   [63:0] reg_2239;
    reg   [63:0] reg_2245;
    reg   [63:0] reg_2250;
    reg   [63:0] reg_2257;
    reg   [63:0] reg_2263;
    reg   [63:0] reg_2269;
    reg   [63:0] reg_2274;
    reg   [63:0] reg_2281;
    wire    ap_CS_fsm_pp0_stage34;
    wire    ap_block_pp0_stage34_11001;
    reg   [63:0] reg_2287;
    reg   [63:0] reg_2293;
    reg   [63:0] reg_2299;
    reg   [63:0] reg_2306;
    reg   [63:0] reg_2313;
    reg   [63:0] reg_2320;
    reg   [63:0] reg_2327;
    reg   [63:0] reg_2333;
    reg   [63:0] reg_2339;
    reg   [63:0] reg_2345;
    reg   [63:0] reg_2350;
    wire    ap_CS_fsm_pp0_stage69;
    wire    ap_block_pp0_stage69_11001;
    reg   [63:0] reg_2356;
    wire    ap_CS_fsm_pp0_stage35;
    wire    ap_block_pp0_stage35_11001;
    reg   [63:0] reg_2361;
    reg   [63:0] reg_2367;
    reg   [63:0] reg_2372;
    reg   [63:0] reg_2378;
    reg   [63:0] reg_2383;
    reg   [63:0] reg_2389;
    reg   [63:0] reg_2396;
    reg   [63:0] reg_2402;
    reg   [63:0] reg_2408;
    reg   [63:0] reg_2414;
    reg   [63:0] reg_2420;
    wire    ap_CS_fsm_pp0_stage70;
    wire    ap_block_pp0_stage70_11001;
    reg   [63:0] reg_2426;
    wire    ap_CS_fsm_pp0_stage36;
    wire    ap_block_pp0_stage36_11001;
    reg   [63:0] reg_2432;
    reg   [63:0] reg_2438;
    reg   [63:0] reg_2445;
    wire   [63:0] grp_fu_1862_p2;
    reg   [63:0] reg_2451;
    wire    ap_CS_fsm_pp0_stage38;
    wire    ap_block_pp0_stage38_11001;
    wire    ap_CS_fsm_pp0_stage45;
    wire    ap_block_pp0_stage45_11001;
    wire    ap_CS_fsm_pp0_stage52;
    wire    ap_block_pp0_stage52_11001;
    wire    ap_CS_fsm_pp0_stage59;
    wire    ap_block_pp0_stage59_11001;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [0:0] icmp_ln263_reg_3394_pp0_iter1_reg;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    wire    ap_CS_fsm_pp0_stage21;
    wire    ap_block_pp0_stage21_11001;
    wire    ap_CS_fsm_pp0_stage22;
    wire    ap_block_pp0_stage22_11001;
    wire   [63:0] grp_fu_1867_p2;
    reg   [63:0] reg_2462;
    wire   [63:0] grp_fu_1872_p2;
    reg   [63:0] reg_2475;
    wire   [63:0] grp_fu_1877_p2;
    reg   [63:0] reg_2488;
    wire   [63:0] grp_fu_1882_p2;
    reg   [63:0] reg_2501;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] grp_fu_1887_p2;
    reg   [63:0] reg_2511;
    wire   [63:0] grp_fu_1892_p2;
    reg   [63:0] reg_2521;
    wire   [63:0] grp_fu_1897_p2;
    reg   [63:0] reg_2530;
    reg   [63:0] reg_2540;
    wire    ap_CS_fsm_pp0_stage39;
    wire    ap_block_pp0_stage39_11001;
    wire    ap_CS_fsm_pp0_stage46;
    wire    ap_block_pp0_stage46_11001;
    wire    ap_CS_fsm_pp0_stage53;
    wire    ap_block_pp0_stage53_11001;
    wire    ap_CS_fsm_pp0_stage15;
    wire    ap_block_pp0_stage15_11001;
    reg   [63:0] reg_2550;
    reg   [63:0] reg_2560;
    reg   [63:0] reg_2570;
    reg   [63:0] reg_2580;
    wire    ap_CS_fsm_pp0_stage40;
    wire    ap_block_pp0_stage40_11001;
    wire    ap_CS_fsm_pp0_stage47;
    wire    ap_block_pp0_stage47_11001;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    reg   [63:0] reg_2589;
    reg   [63:0] reg_2598;
    reg   [63:0] reg_2607;
    wire    ap_CS_fsm_pp0_stage41;
    wire    ap_block_pp0_stage41_11001;
    wire    ap_CS_fsm_pp0_stage48;
    wire    ap_block_pp0_stage48_11001;
    wire    ap_CS_fsm_pp0_stage55;
    wire    ap_block_pp0_stage55_11001;
    wire    ap_CS_fsm_pp0_stage62;
    wire    ap_block_pp0_stage62_11001;
    wire   [63:0] grp_sin_or_cos_double_s_fu_1842_ap_return;
    reg   [63:0] reg_2616;
    wire    ap_CS_fsm_pp0_stage43;
    wire    ap_block_pp0_stage43_11001;
    wire    ap_CS_fsm_pp0_stage44;
    wire    ap_block_pp0_stage44_11001;
    wire    ap_CS_fsm_pp0_stage50;
    wire    ap_block_pp0_stage50_11001;
    wire    ap_CS_fsm_pp0_stage51;
    wire    ap_block_pp0_stage51_11001;
    wire    ap_CS_fsm_pp0_stage56;
    wire    ap_block_pp0_stage56_11001;
    wire    ap_CS_fsm_pp0_stage57;
    wire    ap_block_pp0_stage57_11001;
    reg   [63:0] reg_2626;
    reg   [63:0] reg_2636;
    reg   [63:0] reg_2646;
    reg   [63:0] reg_2657;
    reg   [63:0] reg_2668;
    reg   [63:0] reg_2679;
    reg   [63:0] reg_2689;
    reg   [63:0] reg_2700;
    reg   [63:0] reg_2709;
    reg   [63:0] reg_2720;
    reg   [63:0] reg_2725;
    reg   [63:0] reg_2730;
    wire   [63:0] grp_fu_1902_p2;
    reg   [63:0] reg_2736;
    wire   [63:0] grp_fu_1907_p2;
    reg   [63:0] reg_2742;
    wire   [63:0] grp_fu_1912_p2;
    reg   [63:0] reg_2748;
    wire   [63:0] grp_fu_1917_p2;
    reg   [63:0] reg_2754;
    reg   [2:0] idx_5_reg_3286;
    wire   [0:0] icmp_ln218_fu_2768_p2;
    wire   [63:0] zext_ln218_fu_2774_p1;
    reg   [63:0] zext_ln218_reg_3296;
    reg   [63:0] zext_ln218_reg_3296_pp0_iter1_reg;
    wire   [0:0] icmp_ln263_fu_2795_p2;
    reg   [63:0] l_axis_0_load_reg_3478;
    reg   [63:0] this_TLink_0_0_load_1_reg_3484;
    reg   [63:0] this_TLink_1_0_load_1_reg_3492;
    reg   [63:0] this_TLink_2_0_load_1_reg_3500;
    reg   [63:0] this_TLink_3_0_load_1_reg_3508;
    reg   [63:0] this_TLink_0_1_load_1_reg_3515;
    reg   [63:0] this_TLink_1_1_load_1_reg_3523;
    reg   [63:0] this_TLink_2_1_load_1_reg_3531;
    reg   [63:0] this_TLink_3_1_load_1_reg_3538;
    reg   [63:0] this_TLink_0_2_load_1_reg_3546;
    reg   [63:0] this_TLink_1_2_load_1_reg_3554;
    reg   [63:0] this_TLink_2_2_load_1_reg_3561;
    reg   [63:0] this_TLink_3_2_load_1_reg_3569;
    reg   [63:0] this_TLink_0_3_load_1_reg_3577;
    reg   [63:0] this_TLink_1_3_load_1_reg_3584;
    reg   [63:0] this_TLink_2_3_load_1_reg_3591;
    reg   [63:0] this_TLink_3_3_load_1_reg_3599;
    wire   [0:0] or_ln208_fu_2830_p2;
    reg   [0:0] or_ln208_reg_3607;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire   [0:0] and_ln208_fu_2836_p2;
    reg   [0:0] and_ln208_reg_3612;
    wire   [0:0] icmp_ln208_2_fu_2860_p2;
    reg   [0:0] icmp_ln208_2_reg_3621;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire   [0:0] icmp_ln208_3_fu_2866_p2;
    reg   [0:0] icmp_ln208_3_reg_3626;
    wire   [0:0] and_ln208_1_fu_2876_p2;
    reg   [0:0] and_ln208_1_reg_3631;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    wire   [0:0] icmp_ln208_4_fu_2900_p2;
    reg   [0:0] icmp_ln208_4_reg_3640;
    wire   [0:0] icmp_ln208_5_fu_2906_p2;
    reg   [0:0] icmp_ln208_5_reg_3645;
    wire   [0:0] and_ln208_2_fu_2916_p2;
    reg   [0:0] and_ln208_2_reg_3650;
    wire   [0:0] and_ln208_3_fu_2922_p2;
    reg   [0:0] and_ln208_3_reg_3659;
    wire   [2:0] l_axis_1_addr_1_gep_fu_562_p3;
    wire   [0:0] icmp_ln208_6_fu_2945_p2;
    reg   [0:0] icmp_ln208_6_reg_3668;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    wire   [0:0] icmp_ln208_7_fu_2951_p2;
    reg   [0:0] icmp_ln208_7_reg_3673;
    wire   [0:0] and_ln208_4_fu_2961_p2;
    reg   [0:0] and_ln208_4_reg_3678;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_11001;
    wire   [2:0] l_axis_2_addr_1_gep_fu_738_p3;
    wire   [0:0] icmp_ln208_8_fu_2985_p2;
    reg   [0:0] icmp_ln208_8_reg_3687;
    wire   [0:0] icmp_ln208_9_fu_2991_p2;
    reg   [0:0] icmp_ln208_9_reg_3692;
    wire   [0:0] and_ln208_5_fu_3001_p2;
    reg   [0:0] and_ln208_5_reg_3697;
    wire    ap_CS_fsm_pp0_stage16;
    wire    ap_block_pp0_stage16_11001;
    wire   [2:0] l_axis_1_addr_2_gep_fu_746_p3;
    wire   [2:0] this_q_addr_1_gep_fu_754_p3;
    wire   [0:0] icmp_ln208_10_fu_3025_p2;
    reg   [0:0] icmp_ln208_10_reg_3711;
    wire    ap_CS_fsm_pp0_stage18;
    wire    ap_block_pp0_stage18_11001;
    wire   [0:0] icmp_ln208_11_fu_3031_p2;
    reg   [0:0] icmp_ln208_11_reg_3716;
    wire   [0:0] and_ln208_6_fu_3041_p2;
    reg   [0:0] and_ln208_6_reg_3721;
    wire    ap_CS_fsm_pp0_stage19;
    wire    ap_block_pp0_stage19_11001;
    wire   [2:0] l_axis_2_addr_2_gep_fu_876_p3;
    wire   [0:0] icmp_ln208_12_fu_3065_p2;
    reg   [0:0] icmp_ln208_12_reg_3730;
    wire   [0:0] icmp_ln208_13_fu_3071_p2;
    reg   [0:0] icmp_ln208_13_reg_3735;
    wire   [0:0] and_ln208_7_fu_3081_p2;
    reg   [0:0] and_ln208_7_reg_3740;
    wire   [2:0] this_q_addr_2_gep_fu_884_p3;
    wire   [63:0] zext_ln37_fu_3097_p1;
    reg   [63:0] zext_ln37_reg_3749;
    wire    ap_CS_fsm_pp0_stage24;
    wire    ap_block_pp0_stage24_11001;
    reg   [63:0] this_TCurr_0_0_load_reg_3852;
    reg   [63:0] this_TCurr_0_1_load_reg_3859;
    reg   [63:0] this_TCurr_0_3_load_reg_3870;
    reg   [63:0] this_TCurr_1_0_load_reg_3875;
    reg   [63:0] this_TCurr_1_1_load_reg_3882;
    reg   [63:0] this_TCurr_1_3_load_reg_3894;
    reg   [63:0] this_TCurr_2_0_load_reg_3902;
    reg   [63:0] this_TCurr_2_1_load_reg_3909;
    reg   [63:0] this_TCurr_2_3_load_reg_3921;
    reg   [63:0] this_TCurr_3_0_load_reg_3929;
    reg   [63:0] this_TCurr_3_1_load_reg_3935;
    reg   [63:0] this_TCurr_3_3_load_reg_3945;
    wire   [2:0] this_TJoint_3_0_addr_4_gep_fu_1258_p3;
    wire   [2:0] this_TJoint_3_1_addr_4_gep_fu_1266_p3;
    wire   [2:0] this_TJoint_3_2_addr_4_gep_fu_1274_p3;
    wire   [2:0] this_TJoint_0_3_addr_4_gep_fu_1282_p3;
    wire   [2:0] this_TJoint_1_3_addr_4_gep_fu_1290_p3;
    wire   [2:0] this_TJoint_2_3_addr_4_gep_fu_1298_p3;
    wire   [2:0] this_TJoint_3_3_addr_4_gep_fu_1306_p3;
    reg   [63:0] this_TCurr_0_2_load_reg_3988;
    reg   [63:0] this_TCurr_1_2_load_reg_3994;
    reg   [63:0] this_TCurr_2_2_load_reg_4001;
    reg   [63:0] this_TCurr_3_2_load_reg_4008;
    wire   [2:0] this_TJoint_1_0_addr_4_gep_fu_1369_p3;
    wire   [2:0] this_TJoint_0_1_addr_4_gep_fu_1377_p3;
    wire   [2:0] this_TJoint_1_1_addr_4_gep_fu_1427_p3;
    wire   [2:0] this_TJoint_2_1_addr_4_gep_fu_1452_p3;
    wire   [2:0] this_TJoint_1_2_addr_4_gep_fu_1460_p3;
    wire    ap_CS_fsm_pp0_stage58;
    wire    ap_block_pp0_stage58_11001;
    wire   [2:0] this_TJoint_0_0_addr_4_gep_fu_1518_p3;
    wire   [2:0] this_TJoint_2_2_addr_4_gep_fu_1526_p3;
    wire   [2:0] this_TJoint_2_0_addr_4_gep_fu_1552_p3;
    wire   [2:0] this_TJoint_0_2_addr_4_gep_fu_1560_p3;
    reg   [63:0] mul_i94_2_s_reg_4105;
    reg   [63:0] mul_i94_2_2_1_reg_4110;
    reg   [63:0] mul_i94_1_4_reg_4115;
    reg   [63:0] mul_i94_1_1_2_reg_4120;
    reg   [63:0] mul_i94_1_2_2_reg_4125;
    reg   [63:0] mul_i94_2_4_reg_4130;
    reg   [63:0] mul_i94_2_1_2_reg_4135;
    reg   [63:0] mul_i94_2_2_2_reg_4140;
    reg   [63:0] mul_i94_5_reg_4145;
    reg   [63:0] mul_i94_1158_3_reg_4150;
    reg   [63:0] mul_i94_2165_3_reg_4155;
    reg   [63:0] mul_i94_1_5_reg_4160;
    reg   [63:0] mul_i94_1_1_3_reg_4165;
    reg   [63:0] mul_i94_1_2_3_reg_4170;
    reg   [63:0] mul_i94_1_3_3_reg_4175;
    reg   [63:0] mul_i94_2_5_reg_4180;
    reg   [63:0] mul_i94_2_1_3_reg_4185;
    reg   [63:0] mul_i94_2_2_3_reg_4190;
    reg   [63:0] mul_i94_3_5_reg_4195;
    wire    ap_CS_fsm_pp0_stage71;
    wire    ap_block_pp0_stage71_11001;
    reg   [63:0] mul_i94_3_1_3_reg_4200;
    reg   [63:0] mul_i94_3_2_3_reg_4205;
    reg   [63:0] mul_i94_3_3_3_reg_4210;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    grp_sin_or_cos_double_s_fu_1842_ap_start;
    wire    grp_sin_or_cos_double_s_fu_1842_ap_done;
    wire    grp_sin_or_cos_double_s_fu_1842_ap_idle;
    wire    grp_sin_or_cos_double_s_fu_1842_ap_ready;
    reg   [0:0] grp_sin_or_cos_double_s_fu_1842_do_cos;
    reg    grp_sin_or_cos_double_s_fu_1842_ap_start_reg;
    reg    ap_predicate_op247_call_state12_state11;
    reg    ap_predicate_op255_call_state13_state12;
    reg    ap_predicate_op321_call_state19_state18;
    reg    ap_predicate_op331_call_state20_state19;
    reg    ap_predicate_op425_call_state25_state24;
    reg    ap_predicate_op472_call_state26_state25;
    wire    ap_block_pp0_stage11;
    wire    ap_block_pp0_stage12;
    wire    ap_block_pp0_stage18;
    reg    ap_predicate_pred1771_state19;
    wire    ap_block_pp0_stage19;
    reg    ap_predicate_pred1771_state20;
    wire    ap_block_pp0_stage24;
    reg    ap_predicate_pred1811_state25;
    wire    ap_block_pp0_stage25;
    reg    ap_predicate_pred1811_state26;
    wire    ap_block_pp0_stage13;
    wire    ap_block_pp0_stage20;
    wire    ap_CS_fsm_pp0_stage26;
    wire    ap_block_pp0_stage26;
    wire    ap_CS_fsm_pp0_stage30;
    wire    ap_block_pp0_stage30;
    wire    ap_block_pp0_stage31;
    wire    ap_block_pp0_stage32;
    wire    ap_block_pp0_stage37;
    wire    ap_block_pp0_stage38;
    wire    ap_block_pp0_stage37_11001;
    wire    ap_block_pp0_stage39;
    wire    ap_block_pp0_stage43;
    wire    ap_CS_fsm_pp0_stage42;
    wire    ap_block_pp0_stage42_11001;
    wire    ap_block_pp0_stage44;
    wire    ap_block_pp0_stage45;
    wire    ap_CS_fsm_pp0_stage27;
    wire    ap_block_pp0_stage27;
    wire    ap_block_pp0_stage33;
    wire    ap_block_pp0_stage34;
    wire    ap_block_pp0_stage40;
    wire    ap_block_pp0_stage0;
    wire    ap_block_pp0_stage3;
    wire    ap_block_pp0_stage6;
    wire    ap_block_pp0_stage9;
    wire    ap_block_pp0_stage10;
    wire    ap_block_pp0_stage16;
    wire    ap_block_pp0_stage17;
    wire   [2:0] this_TJoint_0_2_addr_2_gep_fu_790_p3;
    wire   [2:0] this_TJoint_0_3_addr_2_gep_fu_798_p3;
    wire   [2:0] this_TJoint_1_3_addr_2_gep_fu_820_p3;
    wire   [2:0] this_TJoint_2_0_addr_2_gep_fu_828_p3;
    wire   [2:0] this_TJoint_2_3_addr_2_gep_fu_836_p3;
    wire   [2:0] this_TJoint_3_0_addr_2_gep_fu_844_p3;
    wire   [2:0] this_TJoint_3_1_addr_2_gep_fu_852_p3;
    wire   [2:0] this_TJoint_3_2_addr_2_gep_fu_860_p3;
    wire   [2:0] this_TJoint_3_3_addr_2_gep_fu_868_p3;
    wire    ap_block_pp0_stage22;
    wire   [2:0] this_TJoint_0_1_addr_3_gep_fu_892_p3;
    wire    ap_block_pp0_stage23;
    wire   [2:0] this_TJoint_0_3_addr_3_gep_fu_900_p3;
    wire   [2:0] this_TJoint_1_0_addr_3_gep_fu_908_p3;
    wire   [2:0] this_TJoint_1_2_addr_3_gep_fu_930_p3;
    wire   [2:0] this_TJoint_1_3_addr_3_gep_fu_938_p3;
    wire   [2:0] this_TJoint_2_1_addr_3_gep_fu_946_p3;
    wire   [2:0] this_TJoint_2_3_addr_3_gep_fu_954_p3;
    wire   [2:0] this_TJoint_3_0_addr_3_gep_fu_962_p3;
    wire   [2:0] this_TJoint_3_1_addr_3_gep_fu_970_p3;
    wire   [2:0] this_TJoint_3_2_addr_3_gep_fu_978_p3;
    wire   [2:0] this_TJoint_3_3_addr_3_gep_fu_986_p3;
    wire   [2:0] this_TJoint_0_0_addr_1_gep_fu_1321_p3;
    wire   [2:0] this_TJoint_1_1_addr_1_gep_fu_1329_p3;
    wire   [2:0] this_TJoint_0_1_addr_1_gep_fu_1337_p3;
    wire   [2:0] this_TJoint_1_0_addr_1_gep_fu_1345_p3;
    wire    ap_block_pp0_stage46;
    wire   [2:0] this_TJoint_1_1_addr_2_gep_fu_1387_p3;
    wire    ap_block_pp0_stage51;
    reg    ap_predicate_pred1771_state52;
    wire   [2:0] this_TJoint_2_2_addr_2_gep_fu_1395_p3;
    wire    ap_block_pp0_stage52;
    wire   [2:0] this_TJoint_1_2_addr_2_gep_fu_1411_p3;
    reg    ap_predicate_pred1771_state53;
    wire   [2:0] this_TJoint_2_1_addr_2_gep_fu_1419_p3;
    wire    ap_block_pp0_stage53;
    wire   [2:0] this_TJoint_0_0_addr_3_gep_fu_1470_p3;
    wire    ap_block_pp0_stage57;
    reg    ap_predicate_pred1811_state58;
    wire   [2:0] this_TJoint_2_2_addr_3_gep_fu_1478_p3;
    wire    ap_block_pp0_stage58;
    wire   [2:0] this_TJoint_0_2_addr_3_gep_fu_1502_p3;
    reg    ap_predicate_pred1811_state59;
    wire   [2:0] this_TJoint_2_0_addr_3_gep_fu_1510_p3;
    wire    ap_block_pp0_stage59;
    wire    ap_block_pp0_stage61;
    reg   [2:0] idx_fu_202;
    wire   [2:0] add_ln218_fu_3087_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_idx_5;
    wire   [63:0] bitcast_ln251_1_fu_3158_p1;
    wire   [63:0] bitcast_ln237_1_fu_3143_p1;
    wire   [63:0] bitcast_ln221_1_fu_3128_p1;
    reg   [63:0] grp_fu_1862_p0;
    reg   [63:0] grp_fu_1862_p1;
    wire    ap_block_pp0_stage35;
    wire    ap_block_pp0_stage41;
    wire    ap_block_pp0_stage42;
    wire    ap_block_pp0_stage47;
    wire    ap_block_pp0_stage48;
    wire    ap_CS_fsm_pp0_stage49;
    wire    ap_block_pp0_stage49;
    wire    ap_block_pp0_stage54;
    wire    ap_block_pp0_stage55;
    wire    ap_block_pp0_stage56;
    wire    ap_block_pp0_stage62;
    wire    ap_block_pp0_stage67;
    wire    ap_block_pp0_stage68;
    wire    ap_block_pp0_stage69;
    wire    ap_block_pp0_stage1;
    wire    ap_block_pp0_stage2;
    wire    ap_block_pp0_stage8;
    wire    ap_block_pp0_stage15;
    reg   [63:0] grp_fu_1867_p0;
    reg   [63:0] grp_fu_1867_p1;
    reg   [63:0] grp_fu_1872_p0;
    reg   [63:0] grp_fu_1872_p1;
    reg   [63:0] grp_fu_1877_p0;
    reg   [63:0] grp_fu_1877_p1;
    reg   [63:0] grp_fu_1882_p0;
    reg   [63:0] grp_fu_1882_p1;
    reg   [63:0] grp_fu_1887_p0;
    reg   [63:0] grp_fu_1887_p1;
    reg   [63:0] grp_fu_1892_p0;
    reg   [63:0] grp_fu_1892_p1;
    reg   [63:0] grp_fu_1897_p0;
    reg   [63:0] grp_fu_1897_p1;
    reg   [63:0] grp_fu_1902_p0;
    reg   [63:0] grp_fu_1902_p1;
    reg   [63:0] grp_fu_1907_p0;
    reg   [63:0] grp_fu_1907_p1;
    reg   [63:0] grp_fu_1912_p0;
    reg   [63:0] grp_fu_1912_p1;
    reg   [63:0] grp_fu_1917_p0;
    reg   [63:0] grp_fu_1917_p1;
    reg   [63:0] grp_fu_1922_p0;
    reg   [63:0] grp_fu_1922_p1;
    wire    ap_CS_fsm_pp0_stage28;
    wire    ap_block_pp0_stage28;
    wire    ap_CS_fsm_pp0_stage29;
    wire    ap_block_pp0_stage29;
    wire    ap_block_pp0_stage60;
    wire    ap_CS_fsm_pp0_stage63;
    wire    ap_block_pp0_stage63;
    wire    ap_CS_fsm_pp0_stage64;
    wire    ap_block_pp0_stage64;
    wire    ap_CS_fsm_pp0_stage65;
    wire    ap_block_pp0_stage65;
    reg   [63:0] grp_fu_1926_p0;
    reg   [63:0] grp_fu_1926_p1;
    reg   [63:0] grp_fu_1930_p0;
    reg   [63:0] grp_fu_1930_p1;
    reg   [63:0] grp_fu_1934_p0;
    reg   [63:0] grp_fu_1934_p1;
    reg   [63:0] grp_fu_1938_p0;
    reg   [63:0] grp_fu_1938_p1;
    reg   [63:0] grp_fu_1942_p0;
    reg   [63:0] grp_fu_1942_p1;
    reg   [63:0] grp_fu_1946_p0;
    reg   [63:0] grp_fu_1946_p1;
    reg   [63:0] grp_fu_1950_p0;
    reg   [63:0] grp_fu_1950_p1;
    reg   [63:0] grp_fu_1954_p0;
    reg   [63:0] grp_fu_1954_p1;
    reg   [63:0] grp_fu_1958_p0;
    reg   [63:0] grp_fu_1958_p1;
    reg   [63:0] grp_fu_1962_p0;
    reg   [63:0] grp_fu_1962_p1;
    reg   [63:0] grp_fu_1966_p0;
    reg   [63:0] grp_fu_1966_p1;
    reg   [63:0] grp_fu_1970_p0;
    reg   [63:0] grp_fu_1970_p1;
    wire    ap_block_pp0_stage5;
    wire    ap_block_pp0_stage21;
    wire   [63:0] bitcast_ln208_fu_2801_p1;
    wire   [10:0] tmp_271_fu_2804_p4;
    wire   [51:0] trunc_ln208_fu_2814_p1;
    wire   [0:0] icmp_ln208_1_fu_2824_p2;
    wire   [0:0] icmp_ln208_fu_2818_p2;
    wire   [0:0] grp_fu_1970_p2;
    wire   [63:0] bitcast_ln208_1_fu_2842_p1;
    wire   [10:0] tmp_273_fu_2846_p4;
    wire   [51:0] trunc_ln208_1_fu_2856_p1;
    wire   [0:0] or_ln208_1_fu_2872_p2;
    wire   [63:0] bitcast_ln208_2_fu_2882_p1;
    wire   [10:0] tmp_275_fu_2886_p4;
    wire   [51:0] trunc_ln208_2_fu_2896_p1;
    wire   [0:0] or_ln208_2_fu_2912_p2;
    wire   [63:0] bitcast_ln208_3_fu_2927_p1;
    wire   [10:0] tmp_278_fu_2931_p4;
    wire   [51:0] trunc_ln208_3_fu_2941_p1;
    wire   [0:0] or_ln208_3_fu_2957_p2;
    wire   [63:0] bitcast_ln208_4_fu_2967_p1;
    wire   [10:0] tmp_280_fu_2971_p4;
    wire   [51:0] trunc_ln208_4_fu_2981_p1;
    wire   [0:0] or_ln208_4_fu_2997_p2;
    wire   [63:0] bitcast_ln208_5_fu_3007_p1;
    wire   [10:0] tmp_282_fu_3011_p4;
    wire   [51:0] trunc_ln208_5_fu_3021_p1;
    wire   [0:0] or_ln208_5_fu_3037_p2;
    wire   [63:0] bitcast_ln208_6_fu_3047_p1;
    wire   [10:0] tmp_284_fu_3051_p4;
    wire   [51:0] trunc_ln208_6_fu_3061_p1;
    wire   [0:0] or_ln208_6_fu_3077_p2;
    wire   [2:0] add_ln267_fu_3092_p2;
    wire   [63:0] bitcast_ln221_fu_3118_p1;
    wire   [63:0] xor_ln221_fu_3122_p2;
    wire   [63:0] bitcast_ln237_fu_3133_p1;
    wire   [63:0] xor_ln237_fu_3137_p2;
    wire   [63:0] bitcast_ln251_fu_3148_p1;
    wire   [63:0] xor_ln251_fu_3152_p2;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage5_00001;
    wire    ap_block_pp0_stage8_00001;
    wire    ap_block_pp0_stage9_00001;
    wire    ap_block_pp0_stage12_00001;
    reg    ap_predicate_pred3106_state13;
    wire    ap_block_pp0_stage15_00001;
    reg    ap_predicate_pred3117_state16;
    wire    ap_block_pp0_stage18_00001;
    reg    ap_predicate_pred3131_state19;
    wire    ap_block_pp0_stage21_00001;
    reg    ap_predicate_pred3144_state22;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [72:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to1;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_block_pp0_stage13_subdone;
    wire    ap_block_pp0_stage14_subdone;
    wire    ap_block_pp0_stage15_subdone;
    wire    ap_block_pp0_stage16_subdone;
    wire    ap_block_pp0_stage17_subdone;
    wire    ap_block_pp0_stage18_subdone;
    wire    ap_block_pp0_stage19_subdone;
    wire    ap_block_pp0_stage20_subdone;
    wire    ap_block_pp0_stage21_subdone;
    wire    ap_block_pp0_stage22_subdone;
    wire    ap_block_pp0_stage24_subdone;
    wire    ap_block_pp0_stage25_subdone;
    wire    ap_block_pp0_stage26_subdone;
    wire    ap_block_pp0_stage27_subdone;
    wire    ap_block_pp0_stage28_subdone;
    wire    ap_block_pp0_stage29_subdone;
    wire    ap_block_pp0_stage30_subdone;
    wire    ap_block_pp0_stage31_subdone;
    wire    ap_block_pp0_stage32_subdone;
    wire    ap_block_pp0_stage33_subdone;
    wire    ap_block_pp0_stage34_subdone;
    wire    ap_block_pp0_stage35_subdone;
    wire    ap_block_pp0_stage36_subdone;
    wire    ap_block_pp0_stage37_subdone;
    wire    ap_block_pp0_stage38_subdone;
    wire    ap_block_pp0_stage39_subdone;
    wire    ap_block_pp0_stage40_subdone;
    wire    ap_block_pp0_stage41_subdone;
    wire    ap_block_pp0_stage42_subdone;
    wire    ap_block_pp0_stage43_subdone;
    wire    ap_block_pp0_stage44_subdone;
    wire    ap_block_pp0_stage45_subdone;
    wire    ap_block_pp0_stage46_subdone;
    wire    ap_block_pp0_stage47_subdone;
    wire    ap_block_pp0_stage48_subdone;
    wire    ap_block_pp0_stage49_subdone;
    wire    ap_block_pp0_stage50_subdone;
    wire    ap_block_pp0_stage51_subdone;
    wire    ap_block_pp0_stage52_subdone;
    wire    ap_block_pp0_stage53_subdone;
    wire    ap_block_pp0_stage54_subdone;
    wire    ap_block_pp0_stage55_subdone;
    wire    ap_block_pp0_stage56_subdone;
    wire    ap_block_pp0_stage57_subdone;
    wire    ap_block_pp0_stage58_subdone;
    wire    ap_block_pp0_stage59_subdone;
    wire    ap_block_pp0_stage60_subdone;
    wire    ap_block_pp0_stage61_subdone;
    wire    ap_block_pp0_stage62_subdone;
    wire    ap_block_pp0_stage63_subdone;
    wire    ap_block_pp0_stage64_subdone;
    wire    ap_block_pp0_stage65_subdone;
    wire    ap_block_pp0_stage66_subdone;
    wire    ap_block_pp0_stage67_subdone;
    wire    ap_block_pp0_stage68_subdone;
    wire    ap_block_pp0_stage69_subdone;
    wire    ap_block_pp0_stage70_subdone;
    wire    ap_block_pp0_stage71_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    reg    ap_condition_2356;
    reg    ap_condition_3574;
    reg    ap_condition_3579;
    reg    ap_condition_3586;
    reg    ap_condition_3591;
    reg    ap_condition_3597;
    reg    ap_condition_3602;
    reg    ap_condition_3607;
    reg    ap_condition_3612;
    reg    ap_condition_3618;
    reg    ap_condition_3623;
    reg    ap_condition_3629;
    reg    ap_condition_3634;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 73'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 grp_sin_or_cos_double_s_fu_1842_ap_start_reg = 1'b0;
        #0 idx_fu_202 = 3'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_forwardKin_Pipeline_VITIS_LOOP_218_3_l_axis_0_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_axis_0_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_axis_0_address0),
        .ce0(l_axis_0_ce0),
        .q0(l_axis_0_q0)
    );

    main_forwardKin_Pipeline_VITIS_LOOP_218_3_l_axis_1_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_axis_1_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_axis_1_address0),
        .ce0(l_axis_1_ce0),
        .q0(l_axis_1_q0)
    );

    main_forwardKin_Pipeline_VITIS_LOOP_218_3_l_axis_2_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_axis_2_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_axis_2_address0),
        .ce0(l_axis_2_ce0),
        .q0(l_axis_2_q0)
    );

    main_sin_or_cos_double_s grp_sin_or_cos_double_s_fu_1842 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_sin_or_cos_double_s_fu_1842_ap_start),
        .ap_done(grp_sin_or_cos_double_s_fu_1842_ap_done),
        .ap_idle(grp_sin_or_cos_double_s_fu_1842_ap_idle),
        .ap_ready(grp_sin_or_cos_double_s_fu_1842_ap_ready),
        .ap_ce(1'b1),
        .t_in(reg_1987),
        .do_cos(grp_sin_or_cos_double_s_fu_1842_do_cos),
        .ap_return(grp_sin_or_cos_double_s_fu_1842_ap_return)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U375 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1862_p0),
        .din1(grp_fu_1862_p1),
        .ce(1'b1),
        .dout(grp_fu_1862_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U376 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1867_p0),
        .din1(grp_fu_1867_p1),
        .ce(1'b1),
        .dout(grp_fu_1867_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U377 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1872_p0),
        .din1(grp_fu_1872_p1),
        .ce(1'b1),
        .dout(grp_fu_1872_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U378 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1877_p0),
        .din1(grp_fu_1877_p1),
        .ce(1'b1),
        .dout(grp_fu_1877_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U379 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1882_p0),
        .din1(grp_fu_1882_p1),
        .ce(1'b1),
        .dout(grp_fu_1882_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U380 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1887_p0),
        .din1(grp_fu_1887_p1),
        .ce(1'b1),
        .dout(grp_fu_1887_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U381 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1892_p0),
        .din1(grp_fu_1892_p1),
        .ce(1'b1),
        .dout(grp_fu_1892_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U382 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1897_p0),
        .din1(grp_fu_1897_p1),
        .ce(1'b1),
        .dout(grp_fu_1897_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U383 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1902_p0),
        .din1(grp_fu_1902_p1),
        .ce(1'b1),
        .dout(grp_fu_1902_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U384 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1907_p0),
        .din1(grp_fu_1907_p1),
        .ce(1'b1),
        .dout(grp_fu_1907_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U385 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1912_p0),
        .din1(grp_fu_1912_p1),
        .ce(1'b1),
        .dout(grp_fu_1912_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_x_U386 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1917_p0),
        .din1(grp_fu_1917_p1),
        .ce(1'b1),
        .dout(grp_fu_1917_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U387 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1922_p0),
        .din1(grp_fu_1922_p1),
        .ce(1'b1),
        .dout(grp_fu_1922_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U388 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1926_p0),
        .din1(grp_fu_1926_p1),
        .ce(1'b1),
        .dout(grp_fu_1926_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U389 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1930_p0),
        .din1(grp_fu_1930_p1),
        .ce(1'b1),
        .dout(grp_fu_1930_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U390 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1934_p0),
        .din1(grp_fu_1934_p1),
        .ce(1'b1),
        .dout(grp_fu_1934_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U391 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1938_p0),
        .din1(grp_fu_1938_p1),
        .ce(1'b1),
        .dout(grp_fu_1938_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U392 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1942_p0),
        .din1(grp_fu_1942_p1),
        .ce(1'b1),
        .dout(grp_fu_1942_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U393 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1946_p0),
        .din1(grp_fu_1946_p1),
        .ce(1'b1),
        .dout(grp_fu_1946_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U394 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1950_p0),
        .din1(grp_fu_1950_p1),
        .ce(1'b1),
        .dout(grp_fu_1950_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U395 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1954_p0),
        .din1(grp_fu_1954_p1),
        .ce(1'b1),
        .dout(grp_fu_1954_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U396 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1958_p0),
        .din1(grp_fu_1958_p1),
        .ce(1'b1),
        .dout(grp_fu_1958_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U397 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1962_p0),
        .din1(grp_fu_1962_p1),
        .ce(1'b1),
        .dout(grp_fu_1962_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U398 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1966_p0),
        .din1(grp_fu_1966_p1),
        .ce(1'b1),
        .dout(grp_fu_1966_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_U399 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1970_p0),
        .din1(grp_fu_1970_p1),
        .ce(1'b1),
        .opcode(5'd1),
        .dout(grp_fu_1970_p2)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage23),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage23_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage23)) begin
                ap_enable_reg_pp0_iter0_reg <= 1'b0;
            end else if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_subdone))) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage72) & (1'b0 == ap_block_pp0_stage72_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_1842_ap_start_reg <= 1'b0;
        end else begin
            if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (ap_predicate_op247_call_state12_state11 == 1'b1) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (ap_predicate_op321_call_state19_state18 == 1'b1) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11) & (ap_predicate_op255_call_state13_state12 == 1'b1) & (1'b0 == ap_block_pp0_stage11_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (ap_predicate_op472_call_state26_state25 == 1'b1) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18) & (ap_predicate_op331_call_state20_state19 == 1'b1) & (1'b0 == ap_block_pp0_stage18_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (ap_predicate_op425_call_state25_state24 == 1'b1) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
                grp_sin_or_cos_double_s_fu_1842_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_1842_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_1842_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            idx_fu_202 <= 3'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage23_11001))) begin
            idx_fu_202 <= add_ln218_fu_3087_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            and_ln208_1_reg_3631 <= and_ln208_1_fu_2876_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9_11001))) begin
            and_ln208_2_reg_3650 <= and_ln208_2_fu_2916_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001))) begin
            and_ln208_3_reg_3659 <= and_ln208_3_fu_2922_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage13) & (1'b0 == ap_block_pp0_stage13_11001))) begin
            and_ln208_4_reg_3678 <= and_ln208_4_fu_2961_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16_11001))) begin
            and_ln208_5_reg_3697 <= and_ln208_5_fu_3001_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage19) & (1'b0 == ap_block_pp0_stage19_11001))) begin
            and_ln208_6_reg_3721 <= and_ln208_6_fu_3041_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001))) begin
            and_ln208_7_reg_3740 <= and_ln208_7_fu_3081_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            and_ln208_reg_3612 <= and_ln208_fu_2836_p2;
            or_ln208_reg_3607  <= or_ln208_fu_2830_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001))) begin
            ap_predicate_pred1771_state19 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
            ap_predicate_pred3131_state19 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage18) & (1'b0 == ap_block_pp0_stage18_11001))) begin
            ap_predicate_pred1771_state20 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
            icmp_ln208_10_reg_3711 <= icmp_ln208_10_fu_3025_p2;
            icmp_ln208_11_reg_3716 <= icmp_ln208_11_fu_3031_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage50) & (1'b0 == ap_block_pp0_stage50_11001))) begin
            ap_predicate_pred1771_state52 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001))) begin
            ap_predicate_pred1771_state53 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001))) begin
            ap_predicate_pred1811_state25 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
            zext_ln37_reg_3749[2 : 0] <= zext_ln37_fu_3097_p1[2 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001))) begin
            ap_predicate_pred1811_state26 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage56) & (1'b0 == ap_block_pp0_stage56_11001))) begin
            ap_predicate_pred1811_state58 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001))) begin
            ap_predicate_pred1811_state59 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage11) & (1'b0 == ap_block_pp0_stage11_11001))) begin
            ap_predicate_pred3106_state13 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001))) begin
            ap_predicate_pred3117_state16 <= ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage20) & (1'b0 == ap_block_pp0_stage20_11001))) begin
            ap_predicate_pred3144_state22 <= (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001))) begin
            icmp_ln208_12_reg_3730 <= icmp_ln208_12_fu_3065_p2;
            icmp_ln208_13_reg_3735 <= icmp_ln208_13_fu_3071_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5_11001))) begin
            icmp_ln208_2_reg_3621 <= icmp_ln208_2_fu_2860_p2;
            icmp_ln208_3_reg_3626 <= icmp_ln208_3_fu_2866_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001))) begin
            icmp_ln208_4_reg_3640 <= icmp_ln208_4_fu_2900_p2;
            icmp_ln208_5_reg_3645 <= icmp_ln208_5_fu_2906_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage12) & (1'b0 == ap_block_pp0_stage12_11001))) begin
            icmp_ln208_6_reg_3668 <= icmp_ln208_6_fu_2945_p2;
            icmp_ln208_7_reg_3673 <= icmp_ln208_7_fu_2951_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15_11001))) begin
            icmp_ln208_8_reg_3687 <= icmp_ln208_8_fu_2985_p2;
            icmp_ln208_9_reg_3692 <= icmp_ln208_9_fu_2991_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            icmp_ln218_reg_3292 <= icmp_ln218_fu_2768_p2;
            icmp_ln263_reg_3394 <= icmp_ln263_fu_2795_p2;
            icmp_ln263_reg_3394_pp0_iter1_reg <= icmp_ln263_reg_3394;
            idx_5_reg_3286 <= ap_sig_allocacmp_idx_5;
            zext_ln218_reg_3296[2 : 0] <= zext_ln218_fu_2774_p1[2 : 0];
            zext_ln218_reg_3296_pp0_iter1_reg[2 : 0] <= zext_ln218_reg_3296[2 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_axis_0_load_reg_3478 <= l_axis_0_q0;
            this_TLink_0_0_load_1_reg_3484 <= this_TLink_0_0_q0;
            this_TLink_0_1_load_1_reg_3515 <= this_TLink_0_1_q0;
            this_TLink_0_2_load_1_reg_3546 <= this_TLink_0_2_q0;
            this_TLink_0_3_load_1_reg_3577 <= this_TLink_0_3_q0;
            this_TLink_1_0_load_1_reg_3492 <= this_TLink_1_0_q0;
            this_TLink_1_1_load_1_reg_3523 <= this_TLink_1_1_q0;
            this_TLink_1_2_load_1_reg_3554 <= this_TLink_1_2_q0;
            this_TLink_1_3_load_1_reg_3584 <= this_TLink_1_3_q0;
            this_TLink_2_0_load_1_reg_3500 <= this_TLink_2_0_q0;
            this_TLink_2_1_load_1_reg_3531 <= this_TLink_2_1_q0;
            this_TLink_2_2_load_1_reg_3561 <= this_TLink_2_2_q0;
            this_TLink_2_3_load_1_reg_3591 <= this_TLink_2_3_q0;
            this_TLink_3_0_load_1_reg_3508 <= this_TLink_3_0_q0;
            this_TLink_3_1_load_1_reg_3538 <= this_TLink_3_1_q0;
            this_TLink_3_2_load_1_reg_3569 <= this_TLink_3_2_q0;
            this_TLink_3_3_load_1_reg_3599 <= this_TLink_3_3_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage70) & (1'b0 == ap_block_pp0_stage70_11001))) begin
            mul_i94_1158_3_reg_4150 <= grp_fu_1926_p2;
            mul_i94_1_1_3_reg_4165 <= grp_fu_1942_p2;
            mul_i94_1_2_3_reg_4170 <= grp_fu_1946_p2;
            mul_i94_1_3_3_reg_4175 <= grp_fu_1950_p2;
            mul_i94_1_5_reg_4160 <= grp_fu_1938_p2;
            mul_i94_2165_3_reg_4155 <= grp_fu_1930_p2;
            mul_i94_2_1_3_reg_4185 <= grp_fu_1958_p2;
            mul_i94_2_2_3_reg_4190 <= grp_fu_1962_p2;
            mul_i94_2_5_reg_4180 <= grp_fu_1954_p2;
            mul_i94_5_reg_4145 <= grp_fu_1922_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69_11001))) begin
            mul_i94_1_1_2_reg_4120 <= grp_fu_1926_p2;
            mul_i94_1_2_2_reg_4125 <= grp_fu_1930_p2;
            mul_i94_1_4_reg_4115   <= grp_fu_1922_p2;
            mul_i94_2_1_2_reg_4135 <= grp_fu_1942_p2;
            mul_i94_2_2_2_reg_4140 <= grp_fu_1946_p2;
            mul_i94_2_4_reg_4130   <= grp_fu_1938_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (1'b0 == ap_block_pp0_stage68_11001))) begin
            mul_i94_2_2_1_reg_4110 <= grp_fu_1946_p2;
            mul_i94_2_s_reg_4105   <= grp_fu_1938_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage71) & (1'b0 == ap_block_pp0_stage71_11001))) begin
            mul_i94_3_1_3_reg_4200 <= grp_fu_1926_p2;
            mul_i94_3_2_3_reg_4205 <= grp_fu_1930_p2;
            mul_i94_3_3_3_reg_4210 <= grp_fu_1934_p2;
            mul_i94_3_5_reg_4195   <= grp_fu_1922_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11) & (1'b0 == ap_block_pp0_stage11_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001)))) begin
            reg_1977 <= l_axis_1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20) & (1'b0 == ap_block_pp0_stage20_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001)))) begin
            reg_1982 <= l_axis_2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            reg_1987 <= this_q_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage25_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage25) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage25_11001)))) begin
            reg_1992 <= this_TJoint_3_0_q0;
            reg_1999 <= this_TJoint_3_1_q0;
            reg_2006 <= this_TJoint_3_2_q0;
            reg_2013 <= this_TJoint_0_3_q0;
            reg_2025 <= this_TJoint_1_3_q0;
            reg_2035 <= this_TJoint_2_3_q0;
            reg_2045 <= this_TJoint_3_3_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31) & (1'b0 == ap_block_pp0_stage31_11001)))) begin
            reg_2052 <= grp_fu_1922_p2;
            reg_2064 <= grp_fu_1930_p2;
            reg_2077 <= grp_fu_1938_p2;
            reg_2089 <= grp_fu_1946_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31) & (1'b0 == ap_block_pp0_stage31_11001)))) begin
            reg_2058 <= grp_fu_1926_p2;
            reg_2070 <= grp_fu_1934_p2;
            reg_2082 <= grp_fu_1942_p2;
            reg_2095 <= grp_fu_1950_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31) & (1'b0 == ap_block_pp0_stage31_11001)))) begin
            reg_2102 <= grp_fu_1954_p2;
            reg_2108 <= grp_fu_1958_p2;
            reg_2114 <= grp_fu_1962_p2;
            reg_2120 <= grp_fu_1966_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)))) begin
            reg_2126 <= grp_fu_1922_p2;
            reg_2132 <= grp_fu_1926_p2;
            reg_2138 <= grp_fu_1930_p2;
            reg_2145 <= grp_fu_1934_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)))) begin
            reg_2152 <= grp_fu_1938_p2;
            reg_2167 <= grp_fu_1946_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)))) begin
            reg_2159 <= grp_fu_1942_p2;
            reg_2174 <= grp_fu_1950_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage32) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage32_11001)))) begin
            reg_2182 <= grp_fu_1954_p2;
            reg_2189 <= grp_fu_1958_p2;
            reg_2196 <= grp_fu_1962_p2;
            reg_2203 <= grp_fu_1966_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)))) begin
            reg_2209 <= grp_fu_1922_p2;
            reg_2214 <= grp_fu_1926_p2;
            reg_2220 <= grp_fu_1930_p2;
            reg_2233 <= grp_fu_1938_p2;
            reg_2239 <= grp_fu_1942_p2;
            reg_2245 <= grp_fu_1946_p2;
            reg_2257 <= grp_fu_1954_p2;
            reg_2263 <= grp_fu_1958_p2;
            reg_2269 <= grp_fu_1962_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)))) begin
            reg_2225 <= grp_fu_1934_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2250 <= grp_fu_1950_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68_11001)))) begin
            reg_2274 <= grp_fu_1966_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)))) begin
            reg_2281 <= grp_fu_1922_p2;
            reg_2287 <= grp_fu_1926_p2;
            reg_2293 <= grp_fu_1930_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2299 <= grp_fu_1934_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)))) begin
            reg_2306 <= grp_fu_1938_p2;
            reg_2320 <= grp_fu_1946_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage34) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2313 <= grp_fu_1942_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (1'b0 == ap_block_pp0_stage68_11001)))) begin
            reg_2327 <= grp_fu_1950_p2;
            reg_2333 <= grp_fu_1954_p2;
            reg_2339 <= grp_fu_1958_p2;
            reg_2345 <= grp_fu_1962_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34_11001)))) begin
            reg_2350 <= grp_fu_1966_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            reg_2356 <= grp_fu_1922_p2;
            reg_2367 <= grp_fu_1930_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage35) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage35_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)))) begin
            reg_2361 <= grp_fu_1926_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69_11001)))) begin
            reg_2372 <= grp_fu_1934_p2;
            reg_2396 <= grp_fu_1950_p2;
            reg_2402 <= grp_fu_1954_p2;
            reg_2408 <= grp_fu_1958_p2;
            reg_2414 <= grp_fu_1962_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage35) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage35_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2378 <= grp_fu_1938_p2;
            reg_2389 <= grp_fu_1946_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (1'b0 == ap_block_pp0_stage68_11001)))) begin
            reg_2383 <= grp_fu_1942_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage70) & (1'b0 == ap_block_pp0_stage70_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35_11001)))) begin
            reg_2420 <= grp_fu_1966_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage36) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage36_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage66) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage66_11001)))) begin
            reg_2426 <= grp_fu_1922_p2;
            reg_2438 <= grp_fu_1930_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage36) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage36_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2432 <= grp_fu_1926_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36) & (1'b0 == ap_block_pp0_stage36_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage70) & (1'b0 == ap_block_pp0_stage70_11001)))) begin
            reg_2445 <= grp_fu_1934_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 
    == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage52) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage45) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage38) 
    & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage38_11001)))) begin
            reg_2451 <= grp_fu_1862_p2;
            reg_2462 <= grp_fu_1867_p2;
            reg_2475 <= grp_fu_1872_p2;
            reg_2488 <= grp_fu_1877_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage59) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38) & (1'b0 == ap_block_pp0_stage38_11001)))) begin
            reg_2501 <= grp_fu_1882_p2;
            reg_2511 <= grp_fu_1887_p2;
            reg_2521 <= grp_fu_1892_p2;
            reg_2530 <= grp_fu_1897_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 
    == 1'd0) & (1'b0 == ap_block_pp0_stage60_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage39_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage46) 
    & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage39) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage39_11001)))) begin
            reg_2540 <= grp_fu_1862_p2;
            reg_2550 <= grp_fu_1867_p2;
            reg_2560 <= grp_fu_1872_p2;
            reg_2570 <= grp_fu_1877_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 
    == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40_11001)))) begin
            reg_2580 <= grp_fu_1862_p2;
            reg_2589 <= grp_fu_1867_p2;
            reg_2598 <= grp_fu_1872_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) & (1'b0 == ap_block_pp0_stage41_11001)))) begin
            reg_2607 <= grp_fu_1862_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage56) & (1'b0 == ap_block_pp0_stage56_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50) & (1'b0 == ap_block_pp0_stage50_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43) & (1'b0 == ap_block_pp0_stage43_11001)))) begin
            reg_2616 <= grp_sin_or_cos_double_s_fu_1842_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47_11001)))) begin
            reg_2626 <= this_TJoint_1_0_q0;
            reg_2636 <= this_TJoint_0_1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)))) begin
            reg_2646 <= this_TJoint_1_1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54_11001)))) begin
            reg_2657 <= this_TJoint_2_1_q0;
            reg_2668 <= this_TJoint_1_2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)))) begin
            reg_2679 <= this_TJoint_0_0_q0;
            reg_2689 <= this_TJoint_2_2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60_11001)))) begin
            reg_2700 <= this_TJoint_2_0_q0;
            reg_2709 <= this_TJoint_0_2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            reg_2720 <= grp_fu_1877_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67_11001)))) begin
            reg_2725 <= grp_fu_1922_p2;
            reg_2730 <= grp_fu_1930_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001)))) begin
            reg_2736 <= grp_fu_1902_p2;
            reg_2742 <= grp_fu_1907_p2;
            reg_2748 <= grp_fu_1912_p2;
            reg_2754 <= grp_fu_1917_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001))) begin
            this_TCurr_0_0_load_reg_3852 <= this_TCurr_0_0_q0;
            this_TCurr_0_1_load_reg_3859 <= this_TCurr_0_1_q0;
            this_TCurr_0_3_load_reg_3870 <= this_TCurr_0_3_q0;
            this_TCurr_1_0_load_reg_3875 <= this_TCurr_1_0_q0;
            this_TCurr_1_1_load_reg_3882 <= this_TCurr_1_1_q0;
            this_TCurr_1_3_load_reg_3894 <= this_TCurr_1_3_q0;
            this_TCurr_2_0_load_reg_3902 <= this_TCurr_2_0_q0;
            this_TCurr_2_1_load_reg_3909 <= this_TCurr_2_1_q0;
            this_TCurr_2_3_load_reg_3921 <= this_TCurr_2_3_q0;
            this_TCurr_3_0_load_reg_3929 <= this_TCurr_3_0_q0;
            this_TCurr_3_1_load_reg_3935 <= this_TCurr_3_1_q0;
            this_TCurr_3_3_load_reg_3945 <= this_TCurr_3_3_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25_11001))) begin
            this_TCurr_0_2_load_reg_3988 <= this_TCurr_0_2_q0;
            this_TCurr_1_2_load_reg_3994 <= this_TCurr_1_2_q0;
            this_TCurr_2_2_load_reg_4001 <= this_TCurr_2_2_q0;
            this_TCurr_3_2_load_reg_4008 <= this_TCurr_3_2_q0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (icmp_ln218_reg_3292 == 1'd1) & (1'b0 == ap_block_pp0_stage23_subdone))) begin
            ap_condition_exit_pp0_iter0_stage23 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage23 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage23) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage23_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b0)) begin
            ap_idle_pp0_1to1 = 1'b1;
        end else begin
            ap_idle_pp0_1to1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage72) & (1'b0 == ap_block_pp0_stage72_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_idx_5 = 3'd0;
        end else begin
            ap_sig_allocacmp_idx_5 = idx_fu_202;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1862_p0 = reg_2432;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1862_p0 = reg_2730;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)))) begin
            grp_fu_1862_p0 = reg_2426;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1862_p0 = reg_2058;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49) & (1'b0 == ap_block_pp0_stage49)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42) & (1'b0 == ap_block_pp0_stage42)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage56) & (1'b0 == ap_block_pp0_stage56)))) begin
            grp_fu_1862_p0 = reg_2607;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) 
    & (1'b0 == ap_block_pp0_stage41)))) begin
            grp_fu_1862_p0 = reg_2580;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 
    1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1862_p0 = reg_2540;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1862_p0 = reg_2451;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35))) begin
            grp_fu_1862_p0 = reg_2350;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34))) begin
            grp_fu_1862_p0 = reg_2225;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1862_p0 = reg_2126;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1862_p0 = reg_2138;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1862_p0 = reg_2052;
        end else begin
            grp_fu_1862_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
            grp_fu_1862_p1 = mul_i94_2165_3_reg_4155;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1862_p1 = mul_i94_5_reg_4145;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_1862_p1 = reg_2214;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1862_p1 = reg_2299;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1862_p1 = reg_2052;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)))) begin
            grp_fu_1862_p1 = reg_2725;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage56) & (1'b0 == ap_block_pp0_stage56))) begin
            grp_fu_1862_p1 = reg_2445;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1862_p1 = reg_2426;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1862_p1 = reg_2225;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)))) begin
            grp_fu_1862_p1 = reg_2356;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)))) begin
            grp_fu_1862_p1 = reg_2209;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49) & (1'b0 == ap_block_pp0_stage49))) begin
            grp_fu_1862_p1 = reg_2420;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1862_p1 = reg_2361;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)))) begin
            grp_fu_1862_p1 = reg_2138;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1862_p1 = reg_2287;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)))) begin
            grp_fu_1862_p1 = reg_2126;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42) & (1'b0 == ap_block_pp0_stage42))) begin
            grp_fu_1862_p1 = reg_2414;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) & (1'b0 == ap_block_pp0_stage41))) begin
            grp_fu_1862_p1 = reg_2293;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40))) begin
            grp_fu_1862_p1 = reg_2132;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1862_p1 = reg_2220;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1862_p1 = reg_2058;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35) & (1'b0 == ap_block_pp0_stage35)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) 
    & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)))) begin
            grp_fu_1862_p1 = 64'd0;
        end else begin
            grp_fu_1862_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1867_p0 = reg_2299;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1867_p0 = reg_2438;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1867_p0 = reg_2361;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1867_p0 = reg_2070;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) 
    & (1'b0 == ap_block_pp0_stage41)))) begin
            grp_fu_1867_p0 = reg_2589;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 
    1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1867_p0 = reg_2550;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1867_p0 = reg_2462;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)))) begin
            grp_fu_1867_p0 = reg_2250;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1867_p0 = reg_2145;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1867_p0 = reg_2159;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1867_p0 = reg_2064;
        end else begin
            grp_fu_1867_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
            grp_fu_1867_p1 = mul_i94_1_2_3_reg_4170;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1867_p1 = reg_2233;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1867_p1 = mul_i94_1158_3_reg_4150;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1867_p1 = reg_2225;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1867_p1 = mul_i94_1_2_2_reg_4125;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1867_p1 = reg_2730;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_1867_p1 = reg_2239;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1867_p1 = reg_2070;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1867_p1 = reg_2182;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1867_p1 = reg_2064;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1867_p1 = reg_2432;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1867_p1 = reg_2250;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)))) begin
            grp_fu_1867_p1 = reg_2367;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1867_p1 = reg_2281;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1867_p1 = reg_2372;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1867_p1 = reg_2159;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1867_p1 = reg_2306;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1867_p1 = reg_2214;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) & (1'b0 == ap_block_pp0_stage41))) begin
            grp_fu_1867_p1 = reg_2313;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40))) begin
            grp_fu_1867_p1 = reg_2152;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1867_p1 = reg_2245;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1867_p1 = reg_2132;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 
    == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)))) begin
            grp_fu_1867_p1 = 64'd0;
        end else begin
            grp_fu_1867_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1872_p0 = reg_2313;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1872_p0 = reg_2196;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1872_p0 = reg_2306;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1872_p0 = reg_2438;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1872_p0 = reg_2082;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) 
    & (1'b0 == ap_block_pp0_stage41)))) begin
            grp_fu_1872_p0 = reg_2598;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 
    1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1872_p0 = reg_2560;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1872_p0 = reg_2475;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34))) begin
            grp_fu_1872_p0 = reg_2274;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1872_p0 = reg_2167;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1872_p0 = reg_2182;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1872_p0 = reg_2070;
        end else begin
            grp_fu_1872_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
            grp_fu_1872_p1 = mul_i94_2_2_3_reg_4190;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1872_p1 = reg_2257;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1872_p1 = reg_2445;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1872_p1 = reg_2159;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1872_p1 = mul_i94_2_2_2_reg_4140;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_1872_p1 = reg_2263;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1872_p1 = reg_2082;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1872_p1 = mul_i94_2_2_1_reg_4110;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69))) begin
            grp_fu_1872_p1 = reg_2152;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1872_p1 = reg_2138;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1872_p1 = reg_2438;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1872_p1 = reg_2274;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)))) begin
            grp_fu_1872_p1 = reg_2378;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1872_p1 = reg_2233;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1872_p1 = reg_2389;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1872_p1 = reg_2182;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1872_p1 = reg_2327;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)))) begin
            grp_fu_1872_p1 = reg_2145;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41) & (1'b0 == ap_block_pp0_stage41))) begin
            grp_fu_1872_p1 = reg_2383;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40))) begin
            grp_fu_1872_p1 = reg_2174;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1872_p1 = reg_2269;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1872_p1 = reg_2077;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34) & (1'b0 == ap_block_pp0_stage34)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage55)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 
    == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)))) begin
            grp_fu_1872_p1 = 64'd0;
        end else begin
            grp_fu_1872_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68))) begin
            grp_fu_1877_p0 = reg_2250;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1877_p0 = reg_2320;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1877_p0 = reg_2225;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1877_p0 = reg_2720;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1877_p0 = reg_2095;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 
    1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1877_p0 = reg_2570;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1877_p0 = reg_2488;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33))) begin
            grp_fu_1877_p0 = reg_2189;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)))) begin
            grp_fu_1877_p0 = reg_2203;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1877_p0 = reg_2082;
        end else begin
            grp_fu_1877_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
            grp_fu_1877_p1 = reg_2293;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
            grp_fu_1877_p1 = mul_i94_3_2_3_reg_4205;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1877_p1 = reg_2281;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1877_p1 = mul_i94_1_5_reg_4160;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1877_p1 = reg_2174;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1877_p1 = reg_2414;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1877_p1 = reg_2389;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1877_p1 = mul_i94_1_4_reg_4115;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_1877_p1 = reg_2287;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_1877_p1 = reg_2095;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1877_p1 = reg_2089;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1877_p1 = reg_2313;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage69) & (1'b0 == ap_block_pp0_stage69))) begin
            grp_fu_1877_p1 = reg_2167;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1877_p1 = reg_2145;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1877_p1 = reg_2408;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)))) begin
            grp_fu_1877_p1 = reg_2299;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1877_p1 = reg_2203;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage47) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage47))) begin
            grp_fu_1877_p1 = reg_2402;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1877_p1 = reg_2239;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40))) begin
            grp_fu_1877_p1 = reg_2196;
        end else if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage40) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage40)))) begin
            grp_fu_1877_p1 = reg_2345;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39))) begin
            grp_fu_1877_p1 = reg_2152;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage33) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage33)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage67) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 
    == ap_CS_fsm_pp0_stage68) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage68)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1877_p1 = 64'd0;
        end else begin
            grp_fu_1877_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1882_p0 = reg_2306;
        end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1882_p0 = reg_2501;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1882_p0 = reg_2089;
        end else begin
            grp_fu_1882_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1882_p1 = mul_i94_1_1_3_reg_4165;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1882_p1 = mul_i94_1_1_2_reg_4120;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1882_p1 = reg_2389;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1882_p1 = reg_2257;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1882_p1 = reg_2167;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39))) begin
            grp_fu_1882_p1 = reg_2095;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)))) begin
            grp_fu_1882_p1 = 64'd0;
        end else begin
            grp_fu_1882_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1887_p0 = reg_2159;
        end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1887_p0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1887_p0 = reg_2102;
        end else begin
            grp_fu_1887_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1887_p1 = mul_i94_1_3_3_reg_4175;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1887_p1 = reg_2372;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1887_p1 = reg_2189;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1887_p1 = reg_2320;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1887_p1 = reg_2263;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39))) begin
            grp_fu_1887_p1 = reg_2174;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)))) begin
            grp_fu_1887_p1 = 64'd0;
        end else begin
            grp_fu_1887_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1892_p0 = reg_2320;
        end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1892_p0 = reg_2521;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1892_p0 = reg_2108;
        end else begin
            grp_fu_1892_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1892_p1 = mul_i94_2_5_reg_4180;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1892_p1 = mul_i94_2_4_reg_4130;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1892_p1 = mul_i94_2_s_reg_4105;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1892_p1 = reg_2333;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1892_p1 = reg_2189;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39))) begin
            grp_fu_1892_p1 = reg_2114;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)))) begin
            grp_fu_1892_p1 = 64'd0;
        end else begin
            grp_fu_1892_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1897_p0 = reg_2174;
        end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39)))) begin
            grp_fu_1897_p0 = reg_2530;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32))) begin
            grp_fu_1897_p0 = reg_2120;
        end else begin
            grp_fu_1897_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1897_p1 = mul_i94_2_1_3_reg_4185;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1897_p1 = mul_i94_2_1_2_reg_4135;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1897_p1 = reg_2383;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (1'b0 == ap_block_pp0_stage53))) begin
            grp_fu_1897_p1 = reg_2396;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (1'b0 == ap_block_pp0_stage46))) begin
            grp_fu_1897_p1 = reg_2339;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39) & (1'b0 == ap_block_pp0_stage39))) begin
            grp_fu_1897_p1 = reg_2196;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32) & (1'b0 == ap_block_pp0_stage32)))) begin
            grp_fu_1897_p1 = 64'd0;
        end else begin
            grp_fu_1897_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1902_p0 = reg_2736;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1902_p0 = reg_2102;
        end else begin
            grp_fu_1902_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1902_p1 = reg_2420;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1902_p1 = reg_2396;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1902_p1 = reg_2327;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1902_p1 = 64'd0;
        end else begin
            grp_fu_1902_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1907_p0 = reg_2742;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1907_p0 = reg_2108;
        end else begin
            grp_fu_1907_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1907_p1 = mul_i94_3_5_reg_4195;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1907_p1 = reg_2402;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1907_p1 = reg_2333;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1907_p1 = 64'd0;
        end else begin
            grp_fu_1907_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1912_p0 = reg_2748;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1912_p0 = reg_2114;
        end else begin
            grp_fu_1912_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1912_p1 = mul_i94_3_1_3_reg_4200;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1912_p1 = reg_2408;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1912_p1 = reg_2339;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1912_p1 = 64'd0;
        end else begin
            grp_fu_1912_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1917_p0 = reg_2754;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1917_p0 = reg_2120;
        end else begin
            grp_fu_1917_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
            grp_fu_1917_p1 = mul_i94_3_3_3_reg_4210;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
            grp_fu_1917_p1 = reg_2350;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_1917_p1 = reg_2274;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage67) & (1'b0 == ap_block_pp0_stage67))) begin
            grp_fu_1917_p1 = 64'd0;
        end else begin
            grp_fu_1917_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65))) begin
            grp_fu_1922_p0 = reg_2607;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1922_p0 = reg_2580;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1922_p0 = reg_2550;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1922_p0 = reg_2540;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1922_p0 = reg_2462;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1922_p0 = reg_2451;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1922_p0 = this_TLink_0_2_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1922_p0 = this_TLink_0_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1922_p0 = this_TLink_3_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1922_p0 = this_TLink_0_3_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30)))) begin
            grp_fu_1922_p0 = this_TCurr_0_3_load_reg_3870;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)))) begin
            grp_fu_1922_p0 = this_TLink_0_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1922_p0 = this_TCurr_0_2_load_reg_3988;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1922_p0 = this_TCurr_0_0_load_reg_3852;
        end else begin
            grp_fu_1922_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1922_p1 = reg_2700;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)))) begin
            grp_fu_1922_p1 = reg_2679;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1922_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1922_p1 = reg_2646;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1922_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1922_p1 = this_TLink_3_3_load_1_reg_3599;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1922_p1 = this_TLink_3_2_load_1_reg_3569;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1922_p1 = this_TLink_3_1_load_1_reg_3538;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1922_p1 = reg_1992;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1922_p1 = this_TLink_3_0_load_1_reg_3508;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1922_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1922_p1 = this_TLink_2_0_load_1_reg_3500;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1922_p1 = this_TLink_0_0_load_1_reg_3484;
        end else begin
            grp_fu_1922_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65))) begin
            grp_fu_1926_p0 = reg_2607;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1926_p0 = reg_2580;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1926_p0 = reg_2550;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1926_p0 = reg_2540;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1926_p0 = reg_2462;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1926_p0 = this_TLink_0_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1926_p0 = reg_2451;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1926_p0 = this_TLink_1_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1926_p0 = this_TLink_0_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1926_p0 = this_TCurr_1_3_load_reg_3894;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1926_p0 = this_TLink_3_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1926_p0 = this_TLink_0_3_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)))) begin
            grp_fu_1926_p0 = this_TCurr_0_2_load_reg_3988;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1926_p0 = this_TLink_0_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1926_p0 = this_TCurr_0_1_load_reg_3859;
        end else begin
            grp_fu_1926_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1926_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1926_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1926_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1926_p1 = reg_2668;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)))) begin
            grp_fu_1926_p1 = reg_2646;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1926_p1 = reg_2636;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1926_p1 = this_TLink_3_3_load_1_reg_3599;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1926_p1 = this_TLink_2_3_load_1_reg_3591;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1926_p1 = this_TLink_2_2_load_1_reg_3561;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1926_p1 = reg_1999;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1926_p1 = this_TLink_2_1_load_1_reg_3531;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1926_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1926_p1 = this_TLink_1_1_load_1_reg_3523;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1926_p1 = this_TLink_1_0_load_1_reg_3492;
        end else begin
            grp_fu_1926_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65))) begin
            grp_fu_1930_p0 = reg_2607;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1930_p0 = reg_2580;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1930_p0 = reg_2550;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1930_p0 = reg_2540;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1930_p0 = this_TLink_1_0_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)))) begin
            grp_fu_1930_p0 = reg_2451;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1930_p0 = this_TLink_1_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1930_p0 = this_TLink_2_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1930_p0 = this_TLink_1_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1930_p0 = this_TCurr_2_3_load_reg_3921;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1930_p0 = this_TCurr_1_3_load_reg_3894;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1930_p0 = this_TLink_3_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1930_p0 = this_TLink_0_3_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)))) begin
            grp_fu_1930_p0 = this_TCurr_0_1_load_reg_3859;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1930_p0 = this_TLink_0_2_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1930_p0 = this_TCurr_0_0_load_reg_3852;
        end else begin
            grp_fu_1930_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1930_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1930_p1 = reg_2700;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1930_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1930_p1 = reg_2679;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1930_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1930_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1930_p1 = reg_2646;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1930_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1930_p1 = this_TLink_3_3_load_1_reg_3599;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1930_p1 = this_TLink_3_2_load_1_reg_3569;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1930_p1 = this_TLink_1_3_load_1_reg_3584;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1930_p1 = reg_2006;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1930_p1 = this_TLink_1_2_load_1_reg_3554;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1930_p1 = reg_2035;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1930_p1 = this_TLink_0_2_load_1_reg_3546;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1930_p1 = this_TLink_0_1_load_1_reg_3515;
        end else begin
            grp_fu_1930_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65))) begin
            grp_fu_1934_p0 = reg_2607;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1934_p0 = reg_2580;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1934_p0 = reg_2550;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1934_p0 = reg_2540;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1934_p0 = reg_2462;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1934_p0 = this_TLink_1_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1934_p0 = reg_2475;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1934_p0 = this_TLink_1_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1934_p0 = this_TLink_3_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1934_p0 = this_TCurr_3_3_load_reg_3945;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1934_p0 = this_TLink_3_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1934_p0 = this_TCurr_1_3_load_reg_3894;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1934_p0 = this_TLink_0_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1934_p0 = this_TCurr_0_0_load_reg_3852;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1934_p0 = this_TLink_1_0_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)))) begin
            grp_fu_1934_p0 = this_TCurr_1_2_load_reg_3994;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1934_p0 = this_TCurr_1_0_load_reg_3875;
        end else begin
            grp_fu_1934_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1934_p1 = reg_2035;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1934_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1934_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1934_p1 = reg_2679;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1934_p1 = reg_2668;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage54) & (1'b0 == ap_block_pp0_stage54))) begin
            grp_fu_1934_p1 = reg_2646;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1934_p1 = reg_2636;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_1934_p1 = this_TLink_3_3_load_1_reg_3599;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1934_p1 = this_TLink_2_3_load_1_reg_3591;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1934_p1 = this_TLink_3_1_load_1_reg_3538;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage28)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage65) & (1'b0 == ap_block_pp0_stage65)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1934_p1 = reg_2045;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1934_p1 = this_TLink_0_3_load_1_reg_3577;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1934_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1934_p1 = this_TLink_2_0_load_1_reg_3500;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1934_p1 = this_TLink_0_0_load_1_reg_3484;
        end else begin
            grp_fu_1934_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1938_p0 = reg_2589;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1938_p0 = reg_2560;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1938_p0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1938_p0 = reg_2462;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1938_p0 = this_TLink_2_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1938_p0 = reg_2475;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1938_p0 = this_TLink_2_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1938_p0 = this_TLink_2_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1938_p0 = this_TCurr_2_3_load_reg_3921;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1938_p0 = this_TCurr_1_2_load_reg_3994;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1938_p0 = this_TLink_1_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1938_p0 = this_TCurr_1_3_load_reg_3894;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1938_p0 = this_TLink_1_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1938_p0 = this_TCurr_1_1_load_reg_3882;
        end else begin
            grp_fu_1938_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)))) begin
            grp_fu_1938_p1 = reg_2700;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1938_p1 = reg_2679;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1938_p1 = reg_2636;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1938_p1 = reg_2657;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1938_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1938_p1 = this_TLink_3_2_load_1_reg_3569;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1938_p1 = this_TLink_2_2_load_1_reg_3561;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1938_p1 = reg_1992;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1938_p1 = this_TLink_3_0_load_1_reg_3508;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)))) begin
            grp_fu_1938_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1938_p1 = this_TLink_1_1_load_1_reg_3523;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1938_p1 = this_TLink_1_0_load_1_reg_3492;
        end else begin
            grp_fu_1938_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1942_p0 = reg_2589;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1942_p0 = reg_2560;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1942_p0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1942_p0 = reg_2488;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1942_p0 = this_TLink_2_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1942_p0 = reg_2475;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1942_p0 = this_TLink_2_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1942_p0 = this_TLink_2_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1942_p0 = this_TCurr_2_1_load_reg_3909;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1942_p0 = this_TCurr_1_1_load_reg_3882;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1942_p0 = this_TLink_1_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1942_p0 = this_TCurr_1_2_load_reg_3994;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1942_p0 = this_TLink_1_2_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1942_p0 = this_TCurr_1_0_load_reg_3875;
        end else begin
            grp_fu_1942_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1942_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1942_p1 = reg_2646;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1942_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1942_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1942_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1942_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1942_p1 = reg_2668;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1942_p1 = reg_2636;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1942_p1 = this_TLink_1_3_load_1_reg_3584;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1942_p1 = reg_1999;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1942_p1 = this_TLink_2_1_load_1_reg_3531;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1942_p1 = reg_2035;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1942_p1 = this_TLink_0_2_load_1_reg_3546;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1942_p1 = this_TLink_0_1_load_1_reg_3515;
        end else begin
            grp_fu_1942_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1946_p0 = reg_2589;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1946_p0 = reg_2560;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1946_p0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1946_p0 = reg_2488;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1946_p0 = this_TLink_3_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1946_p0 = reg_2501;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55)))) begin
            grp_fu_1946_p0 = this_TLink_3_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1946_p0 = this_TLink_3_1_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1946_p0 = this_TCurr_2_3_load_reg_3921;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1946_p0 = this_TLink_1_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1946_p0 = this_TCurr_1_1_load_reg_3882;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1946_p0 = this_TLink_2_0_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)))) begin
            grp_fu_1946_p0 = this_TCurr_2_2_load_reg_4001;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1946_p0 = this_TCurr_2_0_load_reg_3902;
        end else begin
            grp_fu_1946_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1946_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1946_p1 = reg_2668;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1946_p1 = reg_2700;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1946_p1 = reg_2646;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)))) begin
            grp_fu_1946_p1 = reg_2679;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1946_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48))) begin
            grp_fu_1946_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1946_p1 = this_TLink_2_3_load_1_reg_3591;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1946_p1 = this_TLink_3_1_load_1_reg_3538;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1946_p1 = reg_2006;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1946_p1 = this_TLink_1_2_load_1_reg_3554;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1946_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1946_p1 = this_TLink_2_0_load_1_reg_3500;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1946_p1 = this_TLink_0_0_load_1_reg_3484;
        end else begin
            grp_fu_1946_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1950_p0 = reg_2589;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1950_p0 = reg_2560;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1950_p0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1950_p0 = reg_2475;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1950_p0 = this_TLink_3_2_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1950_p0 = reg_2501;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1950_p0 = this_TLink_3_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1950_p0 = this_TLink_3_0_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1950_p0 = this_TCurr_3_3_load_reg_3945;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1950_p0 = this_TCurr_2_2_load_reg_4001;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1950_p0 = this_TLink_1_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1950_p0 = this_TCurr_1_0_load_reg_3875;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1950_p0 = this_TLink_2_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1950_p0 = this_TCurr_2_1_load_reg_3909;
        end else begin
            grp_fu_1950_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1950_p1 = reg_2035;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61)))) begin
            grp_fu_1950_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1950_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage55) & (1'b0 == ap_block_pp0_stage55))) begin
            grp_fu_1950_p1 = reg_2668;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage60) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48) & (1'b0 == ap_block_pp0_stage48)))) begin
            grp_fu_1950_p1 = reg_2636;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1950_p1 = this_TLink_3_1_load_1_reg_3538;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1950_p1 = this_TLink_2_2_load_1_reg_3561;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1950_p1 = reg_2045;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1950_p1 = this_TLink_0_3_load_1_reg_3577;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62)))) begin
            grp_fu_1950_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1950_p1 = this_TLink_1_1_load_1_reg_3523;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1950_p1 = this_TLink_1_0_load_1_reg_3492;
        end else begin
            grp_fu_1950_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1954_p0 = reg_2598;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1954_p0 = reg_2570;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1954_p0 = reg_2530;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1954_p0 = reg_2488;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1954_p0 = reg_2501;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1954_p0 = this_TCurr_3_2_load_reg_4008;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            grp_fu_1954_p0 = this_TCurr_3_3_load_reg_3945;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1954_p0 = this_TLink_2_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1954_p0 = this_TCurr_2_3_load_reg_3921;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1954_p0 = this_TLink_2_2_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)))) begin
            grp_fu_1954_p0 = this_TCurr_2_0_load_reg_3902;
        end else begin
            grp_fu_1954_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1954_p1 = reg_2700;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1954_p1 = reg_2626;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1954_p1 = reg_2668;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1954_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1954_p1 = this_TLink_2_2_load_1_reg_3561;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1954_p1 = reg_1992;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1954_p1 = this_TLink_3_0_load_1_reg_3508;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1954_p1 = reg_2035;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1954_p1 = this_TLink_0_2_load_1_reg_3546;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1954_p1 = this_TLink_0_1_load_1_reg_3515;
        end else begin
            grp_fu_1954_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1958_p0 = reg_2598;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1958_p0 = reg_2570;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1958_p0 = reg_2530;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1958_p0 = reg_2488;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1958_p0 = reg_2521;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1958_p0 = this_TCurr_3_3_load_reg_3945;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1958_p0 = this_TLink_2_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1958_p0 = this_TCurr_2_2_load_reg_4001;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1958_p0 = this_TLink_3_0_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1958_p0 = this_TCurr_3_2_load_reg_4008;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1958_p0 = this_TCurr_3_0_load_reg_3929;
        end else begin
            grp_fu_1958_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1958_p1 = reg_2657;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1958_p1 = reg_2646;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1958_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1958_p1 = reg_2679;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1958_p1 = this_TLink_3_2_load_1_reg_3569;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1958_p1 = reg_1999;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1958_p1 = this_TLink_2_1_load_1_reg_3531;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1958_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1958_p1 = this_TLink_2_0_load_1_reg_3500;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1958_p1 = this_TLink_0_0_load_1_reg_3484;
        end else begin
            grp_fu_1958_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1962_p0 = reg_2598;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1962_p0 = reg_2570;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1962_p0 = reg_2530;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1962_p0 = reg_2501;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1962_p0 = reg_2521;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1962_p0 = this_TLink_2_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1962_p0 = this_TCurr_2_1_load_reg_3909;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1962_p0 = this_TLink_3_1_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1962_p0 = this_TCurr_3_1_load_reg_3935;
        end else begin
            grp_fu_1962_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1962_p1 = reg_2689;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1962_p1 = reg_2668;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1962_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1962_p1 = reg_2636;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1962_p1 = this_TLink_1_3_load_1_reg_3584;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1962_p1 = reg_2006;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1962_p1 = this_TLink_1_2_load_1_reg_3554;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1962_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1962_p1 = this_TLink_1_1_load_1_reg_3523;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1962_p1 = this_TLink_1_0_load_1_reg_3492;
        end else begin
            grp_fu_1962_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64))) begin
            grp_fu_1966_p0 = reg_2598;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63))) begin
            grp_fu_1966_p0 = reg_2570;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1966_p0 = reg_2530;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61)))) begin
            grp_fu_1966_p0 = reg_2521;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1966_p0 = this_TCurr_3_2_load_reg_4008;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1966_p0 = this_TLink_2_3_load;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27))) begin
            grp_fu_1966_p0 = this_TCurr_2_0_load_reg_3902;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1966_p0 = this_TLink_3_2_load;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1966_p0 = this_TCurr_3_0_load_reg_3929;
        end else begin
            grp_fu_1966_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage62) & (1'b0 == ap_block_pp0_stage62))) begin
            grp_fu_1966_p1 = reg_2025;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            grp_fu_1966_p1 = reg_2709;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage60) & (1'b0 == ap_block_pp0_stage60))) begin
            grp_fu_1966_p1 = reg_2013;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29))) begin
            grp_fu_1966_p1 = this_TLink_2_3_load_1_reg_3591;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage64) & (1'b0 == ap_block_pp0_stage64)))) begin
            grp_fu_1966_p1 = reg_2045;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage27)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28)))) begin
            grp_fu_1966_p1 = this_TLink_0_3_load_1_reg_3577;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage63) & (1'b0 == ap_block_pp0_stage63)))) begin
            grp_fu_1966_p1 = reg_2035;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage26) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage26))) begin
            grp_fu_1966_p1 = this_TLink_0_2_load_1_reg_3546;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25))) begin
            grp_fu_1966_p1 = this_TLink_0_1_load_1_reg_3515;
        end else begin
            grp_fu_1966_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1970_p0 = reg_1982;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18) & (1'b0 == ap_block_pp0_stage18)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (1'b0 == ap_block_pp0_stage12)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5)))) begin
            grp_fu_1970_p0 = reg_1977;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)))) begin
            grp_fu_1970_p0 = l_axis_0_load_reg_3478;
        end else begin
            grp_fu_1970_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
            grp_fu_1970_p1 = 64'd13830554455654793216;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18) & (1'b0 == ap_block_pp0_stage18)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)))) begin
            grp_fu_1970_p1 = 64'd4607182418800017408;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (1'b0 == ap_block_pp0_stage12)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)))) begin
            grp_fu_1970_p1 = 64'd0;
        end else begin
            grp_fu_1970_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25) & (ap_predicate_pred1811_state26 == 1'b1) & (1'b0 == ap_block_pp0_stage25)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19) & (ap_predicate_pred1771_state20 == 1'b1) & (1'b0 == ap_block_pp0_stage19)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage12)))) begin
            grp_sin_or_cos_double_s_fu_1842_do_cos = 1'd0;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage11)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (ap_predicate_pred1811_state25 == 1'b1) & (1'b0 == ap_block_pp0_stage24)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18) & (ap_predicate_pred1771_state19 == 1'b1) & (1'b0 == ap_block_pp0_stage18)))) begin
            grp_sin_or_cos_double_s_fu_1842_do_cos = 1'd1;
        end else begin
            grp_sin_or_cos_double_s_fu_1842_do_cos = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_axis_0_ce0 = 1'b1;
        end else begin
            l_axis_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
                l_axis_1_address0 = l_axis_1_addr_2_gep_fu_746_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                l_axis_1_address0 = l_axis_1_addr_1_gep_fu_562_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
                l_axis_1_address0 = zext_ln218_reg_3296;
            end else begin
                l_axis_1_address0 = 'bx;
            end
        end else begin
            l_axis_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)))) begin
            l_axis_1_ce0 = 1'b1;
        end else begin
            l_axis_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage19) & (1'b0 == ap_block_pp0_stage19))) begin
                l_axis_2_address0 = l_axis_2_addr_2_gep_fu_876_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage13) & (1'b0 == ap_block_pp0_stage13))) begin
                l_axis_2_address0 = l_axis_2_addr_1_gep_fu_738_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
                l_axis_2_address0 = zext_ln218_reg_3296;
            end else begin
                l_axis_2_address0 = 'bx;
            end
        end else begin
            l_axis_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19) & (1'b0 == ap_block_pp0_stage19_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13) & (1'b0 == ap_block_pp0_stage13_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001)))) begin
            l_axis_2_ce0 = 1'b1;
        end else begin
            l_axis_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_0_0_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_0_0_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_0_0_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_0_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_0_0_ce0 = 1'b1;
        end else begin
            this_TCurr_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)))) begin
            this_TCurr_0_0_we0 = 1'b1;
        end else begin
            this_TCurr_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_0_1_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
            this_TCurr_0_1_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_0_1_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_0_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_0_1_ce0 = 1'b1;
        end else begin
            this_TCurr_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
                this_TCurr_0_1_d0 = reg_2462;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TCurr_0_1_d0 = reg_2451;
            end else begin
                this_TCurr_0_1_d0 = 'bx;
            end
        end else begin
            this_TCurr_0_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)))) begin
            this_TCurr_0_1_we0 = 1'b1;
        end else begin
            this_TCurr_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_0_2_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_0_2_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24))) begin
            this_TCurr_0_2_address0 = zext_ln37_reg_3749;
        end else begin
            this_TCurr_0_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001)))) begin
            this_TCurr_0_2_ce0 = 1'b1;
        end else begin
            this_TCurr_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_0_2_we0 = 1'b1;
        end else begin
            this_TCurr_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_0_3_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_0_3_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_0_3_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_0_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_0_3_ce0 = 1'b1;
        end else begin
            this_TCurr_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_0_3_d0 = reg_2475;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_0_3_d0 = reg_2540;
        end else begin
            this_TCurr_0_3_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            this_TCurr_0_3_we0 = 1'b1;
        end else begin
            this_TCurr_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_1_0_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_1_0_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_1_0_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_1_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_1_0_ce0 = 1'b1;
        end else begin
            this_TCurr_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_condition_2356)) begin
            if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1)) begin
                this_TCurr_1_0_d0 = reg_2462;
            end else if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0)) begin
                this_TCurr_1_0_d0 = reg_2488;
            end else begin
                this_TCurr_1_0_d0 = 'bx;
            end
        end else begin
            this_TCurr_1_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)))) begin
            this_TCurr_1_0_we0 = 1'b1;
        end else begin
            this_TCurr_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_1_1_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
            this_TCurr_1_1_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_1_1_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_1_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_1_1_ce0 = 1'b1;
        end else begin
            this_TCurr_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
                this_TCurr_1_1_d0 = reg_2501;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TCurr_1_1_d0 = reg_2462;
            end else begin
                this_TCurr_1_1_d0 = 'bx;
            end
        end else begin
            this_TCurr_1_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)))) begin
            this_TCurr_1_1_we0 = 1'b1;
        end else begin
            this_TCurr_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_1_2_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_1_2_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24))) begin
            this_TCurr_1_2_address0 = zext_ln37_reg_3749;
        end else begin
            this_TCurr_1_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001)))) begin
            this_TCurr_1_2_ce0 = 1'b1;
        end else begin
            this_TCurr_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_1_2_we0 = 1'b1;
        end else begin
            this_TCurr_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_1_3_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_1_3_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_1_3_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_1_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_1_3_ce0 = 1'b1;
        end else begin
            this_TCurr_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_1_3_d0 = reg_2511;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_1_3_d0 = reg_2550;
        end else begin
            this_TCurr_1_3_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            this_TCurr_1_3_we0 = 1'b1;
        end else begin
            this_TCurr_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_2_0_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_2_0_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_2_0_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_2_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_2_0_ce0 = 1'b1;
        end else begin
            this_TCurr_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_condition_2356)) begin
            if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1)) begin
                this_TCurr_2_0_d0 = reg_2475;
            end else if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0)) begin
                this_TCurr_2_0_d0 = reg_2521;
            end else begin
                this_TCurr_2_0_d0 = 'bx;
            end
        end else begin
            this_TCurr_2_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)))) begin
            this_TCurr_2_0_we0 = 1'b1;
        end else begin
            this_TCurr_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_2_1_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
            this_TCurr_2_1_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_2_1_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_2_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_2_1_ce0 = 1'b1;
        end else begin
            this_TCurr_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
                this_TCurr_2_1_d0 = reg_2530;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TCurr_2_1_d0 = reg_2475;
            end else begin
                this_TCurr_2_1_d0 = 'bx;
            end
        end else begin
            this_TCurr_2_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)))) begin
            this_TCurr_2_1_we0 = 1'b1;
        end else begin
            this_TCurr_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_2_2_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_2_2_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24))) begin
            this_TCurr_2_2_address0 = zext_ln37_reg_3749;
        end else begin
            this_TCurr_2_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001)))) begin
            this_TCurr_2_2_ce0 = 1'b1;
        end else begin
            this_TCurr_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_2_2_we0 = 1'b1;
        end else begin
            this_TCurr_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_2_3_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_2_3_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_2_3_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_2_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_2_3_ce0 = 1'b1;
        end else begin
            this_TCurr_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_2_3_d0 = reg_2736;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_2_3_d0 = reg_2560;
        end else begin
            this_TCurr_2_3_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            this_TCurr_2_3_we0 = 1'b1;
        end else begin
            this_TCurr_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_3_0_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_3_0_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_3_0_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_3_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_3_0_ce0 = 1'b1;
        end else begin
            this_TCurr_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_condition_2356)) begin
            if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1)) begin
                this_TCurr_3_0_d0 = reg_2488;
            end else if ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0)) begin
                this_TCurr_3_0_d0 = reg_2742;
            end else begin
                this_TCurr_3_0_d0 = 'bx;
            end
        end else begin
            this_TCurr_3_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)))) begin
            this_TCurr_3_0_we0 = 1'b1;
        end else begin
            this_TCurr_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_3_1_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
            this_TCurr_3_1_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_3_1_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_3_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_3_1_ce0 = 1'b1;
        end else begin
            this_TCurr_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
                this_TCurr_3_1_d0 = reg_2748;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TCurr_3_1_d0 = reg_2488;
            end else begin
                this_TCurr_3_1_d0 = 'bx;
            end
        end else begin
            this_TCurr_3_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)))) begin
            this_TCurr_3_1_we0 = 1'b1;
        end else begin
            this_TCurr_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_3_2_address0 = 64'd0;
        end else if (((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_3_2_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24))) begin
            this_TCurr_3_2_address0 = zext_ln37_reg_3749;
        end else begin
            this_TCurr_3_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001)))) begin
            this_TCurr_3_2_ce0 = 1'b1;
        end else begin
            this_TCurr_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)) | ((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_3_2_we0 = 1'b1;
        end else begin
            this_TCurr_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_3_3_address0 = zext_ln218_reg_3296_pp0_iter1_reg;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_3_3_address0 = 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TCurr_3_3_address0 = zext_ln37_fu_3097_p1;
        end else begin
            this_TCurr_3_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TCurr_3_3_ce0 = 1'b1;
        end else begin
            this_TCurr_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
            this_TCurr_3_3_d0 = reg_2754;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (1'b0 == ap_block_pp0_stage61))) begin
            this_TCurr_3_3_d0 = reg_2570;
        end else begin
            this_TCurr_3_3_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((icmp_ln263_reg_3394_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage61) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage61_11001)))) begin
            this_TCurr_3_3_we0 = 1'b1;
        end else begin
            this_TCurr_3_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3579)) begin
                this_TJoint_0_0_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3574)) begin
                this_TJoint_0_0_address0 = this_TJoint_0_0_addr_4_gep_fu_1518_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57))) begin
                this_TJoint_0_0_address0 = this_TJoint_0_0_addr_3_gep_fu_1470_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44))) begin
                this_TJoint_0_0_address0 = this_TJoint_0_0_addr_1_gep_fu_1321_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_0_0_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_0_0_address0 = 'bx;
            end
        end else begin
            this_TJoint_0_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44_11001)))) begin
            this_TJoint_0_0_ce0 = 1'b1;
        end else begin
            this_TJoint_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44)))) begin
            this_TJoint_0_0_d0 = reg_2616;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
            this_TJoint_0_0_d0 = 64'd4607182418800017408;
        end else begin
            this_TJoint_0_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1811_state58 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage44_11001)))) begin
            this_TJoint_0_0_we0 = 1'b1;
        end else begin
            this_TJoint_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3591)) begin
                this_TJoint_0_1_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3586)) begin
                this_TJoint_0_1_address0 = this_TJoint_0_1_addr_4_gep_fu_1377_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45))) begin
                this_TJoint_0_1_address0 = this_TJoint_0_1_addr_1_gep_fu_1337_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_0_1_address0 = this_TJoint_0_1_addr_3_gep_fu_892_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_0_1_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_0_1_address0 = 'bx;
            end
        end else begin
            this_TJoint_0_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_0_1_ce0 = 1'b1;
        end else begin
            this_TJoint_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45))) begin
            this_TJoint_0_1_d0 = bitcast_ln221_1_fu_3128_p1;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23)))) begin
            this_TJoint_0_1_d0 = 64'd0;
        end else begin
            this_TJoint_0_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_0_1_we0 = 1'b1;
        end else begin
            this_TJoint_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3602)) begin
                this_TJoint_0_2_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3597)) begin
                this_TJoint_0_2_address0 = this_TJoint_0_2_addr_4_gep_fu_1560_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58))) begin
                this_TJoint_0_2_address0 = this_TJoint_0_2_addr_3_gep_fu_1502_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_0_2_address0 = this_TJoint_0_2_addr_2_gep_fu_790_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_0_2_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_0_2_address0 = 'bx;
            end
        end else begin
            this_TJoint_0_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58_11001)))) begin
            this_TJoint_0_2_ce0 = 1'b1;
        end else begin
            this_TJoint_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58))) begin
            this_TJoint_0_2_d0 = reg_2616;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17)))) begin
            this_TJoint_0_2_d0 = 64'd0;
        end else begin
            this_TJoint_0_2_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1811_state59 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58_11001)))) begin
            this_TJoint_0_2_we0 = 1'b1;
        end else begin
            this_TJoint_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_0_3_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_0_3_address0 = this_TJoint_0_3_addr_4_gep_fu_1282_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_0_3_address0 = this_TJoint_0_3_addr_3_gep_fu_900_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_0_3_address0 = this_TJoint_0_3_addr_2_gep_fu_798_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_0_3_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_0_3_address0 = 'bx;
            end
        end else begin
            this_TJoint_0_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_0_3_ce0 = 1'b1;
        end else begin
            this_TJoint_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_0_3_we0 = 1'b1;
        end else begin
            this_TJoint_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3591)) begin
                this_TJoint_1_0_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3586)) begin
                this_TJoint_1_0_address0 = this_TJoint_1_0_addr_4_gep_fu_1369_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45))) begin
                this_TJoint_1_0_address0 = this_TJoint_1_0_addr_1_gep_fu_1345_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_1_0_address0 = this_TJoint_1_0_addr_3_gep_fu_908_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_1_0_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_1_0_address0 = 'bx;
            end
        end else begin
            this_TJoint_1_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_1_0_ce0 = 1'b1;
        end else begin
            this_TJoint_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'b0 == ap_block_pp0_stage45))) begin
            this_TJoint_1_0_d0 = reg_2616;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23)))) begin
            this_TJoint_1_0_d0 = 64'd0;
        end else begin
            this_TJoint_1_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage45_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_1_0_we0 = 1'b1;
        end else begin
            this_TJoint_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3623)) begin
                this_TJoint_1_1_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3618)) begin
                this_TJoint_1_1_address0 = this_TJoint_1_1_addr_4_gep_fu_1427_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51))) begin
                this_TJoint_1_1_address0 = this_TJoint_1_1_addr_2_gep_fu_1387_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44))) begin
                this_TJoint_1_1_address0 = this_TJoint_1_1_addr_1_gep_fu_1329_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_1_1_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_1_1_address0 = 'bx;
            end
        end else begin
            this_TJoint_1_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage52) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_1_1_ce0 = 1'b1;
        end else begin
            this_TJoint_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'b0 == ap_block_pp0_stage44)))) begin
            this_TJoint_1_1_d0 = reg_2616;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
            this_TJoint_1_1_d0 = 64'd4607182418800017408;
        end else begin
            this_TJoint_1_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1771_state52 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage44_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) 
    & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_1_1_we0 = 1'b1;
        end else begin
            this_TJoint_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3634)) begin
                this_TJoint_1_2_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3629)) begin
                this_TJoint_1_2_address0 = this_TJoint_1_2_addr_4_gep_fu_1460_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52))) begin
                this_TJoint_1_2_address0 = this_TJoint_1_2_addr_2_gep_fu_1411_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_1_2_address0 = this_TJoint_1_2_addr_3_gep_fu_930_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_1_2_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_1_2_address0 = 'bx;
            end
        end else begin
            this_TJoint_1_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_1_2_ce0 = 1'b1;
        end else begin
            this_TJoint_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52))) begin
            this_TJoint_1_2_d0 = reg_2616;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23)))) begin
            this_TJoint_1_2_d0 = 64'd0;
        end else begin
            this_TJoint_1_2_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1771_state53 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) 
    & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_1_2_we0 = 1'b1;
        end else begin
            this_TJoint_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_1_3_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_1_3_address0 = this_TJoint_1_3_addr_4_gep_fu_1290_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_1_3_address0 = this_TJoint_1_3_addr_3_gep_fu_938_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_1_3_address0 = this_TJoint_1_3_addr_2_gep_fu_820_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_1_3_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_1_3_address0 = 'bx;
            end
        end else begin
            this_TJoint_1_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_1_3_ce0 = 1'b1;
        end else begin
            this_TJoint_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_1_3_we0 = 1'b1;
        end else begin
            this_TJoint_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3602)) begin
                this_TJoint_2_0_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3597)) begin
                this_TJoint_2_0_address0 = this_TJoint_2_0_addr_4_gep_fu_1552_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58))) begin
                this_TJoint_2_0_address0 = this_TJoint_2_0_addr_3_gep_fu_1510_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_2_0_address0 = this_TJoint_2_0_addr_2_gep_fu_828_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_2_0_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_2_0_address0 = 'bx;
            end
        end else begin
            this_TJoint_2_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58_11001)))) begin
            this_TJoint_2_0_ce0 = 1'b1;
        end else begin
            this_TJoint_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58))) begin
            this_TJoint_2_0_d0 = bitcast_ln251_1_fu_3158_p1;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17)))) begin
            this_TJoint_2_0_d0 = 64'd0;
        end else begin
            this_TJoint_2_0_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1811_state59 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (1'b0 == ap_block_pp0_stage58_11001)))) begin
            this_TJoint_2_0_we0 = 1'b1;
        end else begin
            this_TJoint_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3634)) begin
                this_TJoint_2_1_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3629)) begin
                this_TJoint_2_1_address0 = this_TJoint_2_1_addr_4_gep_fu_1452_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52))) begin
                this_TJoint_2_1_address0 = this_TJoint_2_1_addr_2_gep_fu_1419_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_2_1_address0 = this_TJoint_2_1_addr_3_gep_fu_946_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_2_1_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_2_1_address0 = 'bx;
            end
        end else begin
            this_TJoint_2_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_2_1_ce0 = 1'b1;
        end else begin
            this_TJoint_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52))) begin
            this_TJoint_2_1_d0 = bitcast_ln237_1_fu_3143_p1;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23)))) begin
            this_TJoint_2_1_d0 = 64'd0;
        end else begin
            this_TJoint_2_1_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1771_state53 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (1'b0 == ap_block_pp0_stage52_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) 
    & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_2_1_we0 = 1'b1;
        end else begin
            this_TJoint_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3579)) begin
                this_TJoint_2_2_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3574)) begin
                this_TJoint_2_2_address0 = this_TJoint_2_2_addr_4_gep_fu_1526_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57))) begin
                this_TJoint_2_2_address0 = this_TJoint_2_2_addr_3_gep_fu_1478_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51))) begin
                this_TJoint_2_2_address0 = this_TJoint_2_2_addr_2_gep_fu_1395_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_2_2_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_2_2_address0 = 'bx;
            end
        end else begin
            this_TJoint_2_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001)))) begin
            this_TJoint_2_2_ce0 = 1'b1;
        end else begin
            this_TJoint_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51)))) begin
            this_TJoint_2_2_d0 = reg_2616;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
            this_TJoint_2_2_d0 = 64'd4607182418800017408;
        end else begin
            this_TJoint_2_2_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1811_state58 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage57) & (1'b0 == ap_block_pp0_stage57_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_predicate_pred1771_state52 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51) & (1'b0 == ap_block_pp0_stage51_11001)))) begin
            this_TJoint_2_2_we0 = 1'b1;
        end else begin
            this_TJoint_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_2_3_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_2_3_address0 = this_TJoint_2_3_addr_4_gep_fu_1298_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_2_3_address0 = this_TJoint_2_3_addr_3_gep_fu_954_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_2_3_address0 = this_TJoint_2_3_addr_2_gep_fu_836_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_2_3_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_2_3_address0 = 'bx;
            end
        end else begin
            this_TJoint_2_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_2_3_ce0 = 1'b1;
        end else begin
            this_TJoint_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_2_3_we0 = 1'b1;
        end else begin
            this_TJoint_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_3_0_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_3_0_address0 = this_TJoint_3_0_addr_4_gep_fu_1258_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_3_0_address0 = this_TJoint_3_0_addr_3_gep_fu_962_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_3_0_address0 = this_TJoint_3_0_addr_2_gep_fu_844_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_3_0_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_3_0_address0 = 'bx;
            end
        end else begin
            this_TJoint_3_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_3_0_ce0 = 1'b1;
        end else begin
            this_TJoint_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_3_0_we0 = 1'b1;
        end else begin
            this_TJoint_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_3_1_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_3_1_address0 = this_TJoint_3_1_addr_4_gep_fu_1266_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_3_1_address0 = this_TJoint_3_1_addr_3_gep_fu_970_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_3_1_address0 = this_TJoint_3_1_addr_2_gep_fu_852_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_3_1_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_3_1_address0 = 'bx;
            end
        end else begin
            this_TJoint_3_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_3_1_ce0 = 1'b1;
        end else begin
            this_TJoint_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_3_1_we0 = 1'b1;
        end else begin
            this_TJoint_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_3_2_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_3_2_address0 = this_TJoint_3_2_addr_4_gep_fu_1274_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_3_2_address0 = this_TJoint_3_2_addr_3_gep_fu_978_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_3_2_address0 = this_TJoint_3_2_addr_2_gep_fu_860_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_3_2_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_3_2_address0 = 'bx;
            end
        end else begin
            this_TJoint_3_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_3_2_ce0 = 1'b1;
        end else begin
            this_TJoint_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_3_2_we0 = 1'b1;
        end else begin
            this_TJoint_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if ((1'b1 == ap_condition_3612)) begin
                this_TJoint_3_3_address0 = 64'd0;
            end else if ((1'b1 == ap_condition_3607)) begin
                this_TJoint_3_3_address0 = this_TJoint_3_3_addr_4_gep_fu_1306_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23))) begin
                this_TJoint_3_3_address0 = this_TJoint_3_3_addr_3_gep_fu_986_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17))) begin
                this_TJoint_3_3_address0 = this_TJoint_3_3_addr_2_gep_fu_868_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10))) begin
                this_TJoint_3_3_address0 = zext_ln218_reg_3296;
            end else begin
                this_TJoint_3_3_address0 = 'bx;
            end
        end else begin
            this_TJoint_3_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001)))) begin
            this_TJoint_3_3_ce0 = 1'b1;
        end else begin
            this_TJoint_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10) & (1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage10_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17) & (1'b0 == ap_block_pp0_stage17_11001) & ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)))) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001) & (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) 
    & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 
    == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)))))) begin
            this_TJoint_3_3_we0 = 1'b1;
        end else begin
            this_TJoint_3_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_0_0_ce0 = 1'b1;
        end else begin
            this_TLink_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_0_1_ce0 = 1'b1;
        end else begin
            this_TLink_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_0_2_ce0 = 1'b1;
        end else begin
            this_TLink_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_0_3_ce0 = 1'b1;
        end else begin
            this_TLink_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_1_0_ce0 = 1'b1;
        end else begin
            this_TLink_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_1_1_ce0 = 1'b1;
        end else begin
            this_TLink_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_1_2_ce0 = 1'b1;
        end else begin
            this_TLink_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_1_3_ce0 = 1'b1;
        end else begin
            this_TLink_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_2_0_ce0 = 1'b1;
        end else begin
            this_TLink_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_2_1_ce0 = 1'b1;
        end else begin
            this_TLink_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_2_2_ce0 = 1'b1;
        end else begin
            this_TLink_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_2_3_ce0 = 1'b1;
        end else begin
            this_TLink_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_3_0_ce0 = 1'b1;
        end else begin
            this_TLink_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_3_1_ce0 = 1'b1;
        end else begin
            this_TLink_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_3_2_ce0 = 1'b1;
        end else begin
            this_TLink_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            this_TLink_3_3_ce0 = 1'b1;
        end else begin
            this_TLink_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22))) begin
                this_q_address0 = this_q_addr_2_gep_fu_884_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16))) begin
                this_q_address0 = this_q_addr_1_gep_fu_754_p3;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9))) begin
                this_q_address0 = zext_ln218_reg_3296;
            end else begin
                this_q_address0 = 'bx;
            end
        end else begin
            this_q_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9) & (1'b0 == ap_block_pp0_stage9_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16) & (1'b0 == ap_block_pp0_stage16_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001)))) begin
            this_q_ce0 = 1'b1;
        end else begin
            this_q_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to1 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            ap_ST_fsm_pp0_stage14: begin
                if ((1'b0 == ap_block_pp0_stage14_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end
            end
            ap_ST_fsm_pp0_stage15: begin
                if ((1'b0 == ap_block_pp0_stage15_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end
            end
            ap_ST_fsm_pp0_stage16: begin
                if ((1'b0 == ap_block_pp0_stage16_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end
            end
            ap_ST_fsm_pp0_stage17: begin
                if ((1'b0 == ap_block_pp0_stage17_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end
            end
            ap_ST_fsm_pp0_stage18: begin
                if ((1'b0 == ap_block_pp0_stage18_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end
            end
            ap_ST_fsm_pp0_stage19: begin
                if ((1'b0 == ap_block_pp0_stage19_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end
            end
            ap_ST_fsm_pp0_stage20: begin
                if ((1'b0 == ap_block_pp0_stage20_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end
            end
            ap_ST_fsm_pp0_stage21: begin
                if ((1'b0 == ap_block_pp0_stage21_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end
            end
            ap_ST_fsm_pp0_stage22: begin
                if ((1'b0 == ap_block_pp0_stage22_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end
            end
            ap_ST_fsm_pp0_stage23: begin
                if ((1'b1 == ap_condition_exit_pp0_iter0_stage23)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage23_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end
            end
            ap_ST_fsm_pp0_stage24: begin
                if ((1'b0 == ap_block_pp0_stage24_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end
            end
            ap_ST_fsm_pp0_stage25: begin
                if ((1'b0 == ap_block_pp0_stage25_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end
            end
            ap_ST_fsm_pp0_stage26: begin
                if ((1'b0 == ap_block_pp0_stage26_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end
            end
            ap_ST_fsm_pp0_stage27: begin
                if ((1'b0 == ap_block_pp0_stage27_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end
            end
            ap_ST_fsm_pp0_stage28: begin
                if ((1'b0 == ap_block_pp0_stage28_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end
            end
            ap_ST_fsm_pp0_stage29: begin
                if ((1'b0 == ap_block_pp0_stage29_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end
            end
            ap_ST_fsm_pp0_stage30: begin
                if ((1'b0 == ap_block_pp0_stage30_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end
            end
            ap_ST_fsm_pp0_stage31: begin
                if ((1'b0 == ap_block_pp0_stage31_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end
            end
            ap_ST_fsm_pp0_stage32: begin
                if ((1'b0 == ap_block_pp0_stage32_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end
            end
            ap_ST_fsm_pp0_stage33: begin
                if ((1'b0 == ap_block_pp0_stage33_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end
            end
            ap_ST_fsm_pp0_stage34: begin
                if ((1'b0 == ap_block_pp0_stage34_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end
            end
            ap_ST_fsm_pp0_stage35: begin
                if ((1'b0 == ap_block_pp0_stage35_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end
            end
            ap_ST_fsm_pp0_stage36: begin
                if ((1'b0 == ap_block_pp0_stage36_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end
            end
            ap_ST_fsm_pp0_stage37: begin
                if ((1'b0 == ap_block_pp0_stage37_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end
            end
            ap_ST_fsm_pp0_stage38: begin
                if ((1'b0 == ap_block_pp0_stage38_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end
            end
            ap_ST_fsm_pp0_stage39: begin
                if ((1'b0 == ap_block_pp0_stage39_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end
            end
            ap_ST_fsm_pp0_stage40: begin
                if ((1'b0 == ap_block_pp0_stage40_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end
            end
            ap_ST_fsm_pp0_stage41: begin
                if ((1'b0 == ap_block_pp0_stage41_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end
            end
            ap_ST_fsm_pp0_stage42: begin
                if ((1'b0 == ap_block_pp0_stage42_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end
            end
            ap_ST_fsm_pp0_stage43: begin
                if ((1'b0 == ap_block_pp0_stage43_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end
            end
            ap_ST_fsm_pp0_stage44: begin
                if ((1'b0 == ap_block_pp0_stage44_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end
            end
            ap_ST_fsm_pp0_stage45: begin
                if ((1'b0 == ap_block_pp0_stage45_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end
            end
            ap_ST_fsm_pp0_stage46: begin
                if ((1'b0 == ap_block_pp0_stage46_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end
            end
            ap_ST_fsm_pp0_stage47: begin
                if ((1'b0 == ap_block_pp0_stage47_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end
            end
            ap_ST_fsm_pp0_stage48: begin
                if ((1'b0 == ap_block_pp0_stage48_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end
            end
            ap_ST_fsm_pp0_stage49: begin
                if ((1'b0 == ap_block_pp0_stage49_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end
            end
            ap_ST_fsm_pp0_stage50: begin
                if ((1'b0 == ap_block_pp0_stage50_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end
            end
            ap_ST_fsm_pp0_stage51: begin
                if ((1'b0 == ap_block_pp0_stage51_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end
            end
            ap_ST_fsm_pp0_stage52: begin
                if ((1'b0 == ap_block_pp0_stage52_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end
            end
            ap_ST_fsm_pp0_stage53: begin
                if ((1'b0 == ap_block_pp0_stage53_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end
            end
            ap_ST_fsm_pp0_stage54: begin
                if ((1'b0 == ap_block_pp0_stage54_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end
            end
            ap_ST_fsm_pp0_stage55: begin
                if ((1'b0 == ap_block_pp0_stage55_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end
            end
            ap_ST_fsm_pp0_stage56: begin
                if ((1'b0 == ap_block_pp0_stage56_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end
            end
            ap_ST_fsm_pp0_stage57: begin
                if ((1'b0 == ap_block_pp0_stage57_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end
            end
            ap_ST_fsm_pp0_stage58: begin
                if ((1'b0 == ap_block_pp0_stage58_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end
            end
            ap_ST_fsm_pp0_stage59: begin
                if ((1'b0 == ap_block_pp0_stage59_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end
            end
            ap_ST_fsm_pp0_stage60: begin
                if ((1'b0 == ap_block_pp0_stage60_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end
            end
            ap_ST_fsm_pp0_stage61: begin
                if ((1'b0 == ap_block_pp0_stage61_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end
            end
            ap_ST_fsm_pp0_stage62: begin
                if ((1'b0 == ap_block_pp0_stage62_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end
            end
            ap_ST_fsm_pp0_stage63: begin
                if ((1'b0 == ap_block_pp0_stage63_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end
            end
            ap_ST_fsm_pp0_stage64: begin
                if ((1'b0 == ap_block_pp0_stage64_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end
            end
            ap_ST_fsm_pp0_stage65: begin
                if ((1'b0 == ap_block_pp0_stage65_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end
            end
            ap_ST_fsm_pp0_stage66: begin
                if ((1'b0 == ap_block_pp0_stage66_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end
            end
            ap_ST_fsm_pp0_stage67: begin
                if ((1'b0 == ap_block_pp0_stage67_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end
            end
            ap_ST_fsm_pp0_stage68: begin
                if ((1'b0 == ap_block_pp0_stage68_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage69;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end
            end
            ap_ST_fsm_pp0_stage69: begin
                if ((1'b0 == ap_block_pp0_stage69_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage70;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage69;
                end
            end
            ap_ST_fsm_pp0_stage70: begin
                if ((1'b0 == ap_block_pp0_stage70_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage71;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage70;
                end
            end
            ap_ST_fsm_pp0_stage71: begin
                if ((1'b0 == ap_block_pp0_stage71_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage72;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage71;
                end
            end
            ap_ST_fsm_pp0_stage72: begin
                if ((1'b0 == ap_block_pp0_stage72_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage72;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln218_fu_3087_p2 = (idx_5_reg_3286 + 3'd1);

    assign add_ln267_fu_3092_p2 = ($signed(idx_5_reg_3286) + $signed(3'd7));

    assign and_ln208_1_fu_2876_p2 = (or_ln208_1_fu_2872_p2 & grp_fu_1970_p2);

    assign and_ln208_2_fu_2916_p2 = (or_ln208_2_fu_2912_p2 & grp_fu_1970_p2);

    assign and_ln208_3_fu_2922_p2 = (or_ln208_reg_3607 & grp_fu_1970_p2);

    assign and_ln208_4_fu_2961_p2 = (or_ln208_3_fu_2957_p2 & grp_fu_1970_p2);

    assign and_ln208_5_fu_3001_p2 = (or_ln208_4_fu_2997_p2 & grp_fu_1970_p2);

    assign and_ln208_6_fu_3041_p2 = (or_ln208_5_fu_3037_p2 & grp_fu_1970_p2);

    assign and_ln208_7_fu_3081_p2 = (or_ln208_6_fu_3077_p2 & grp_fu_1970_p2);

    assign and_ln208_fu_2836_p2 = (or_ln208_fu_2830_p2 & grp_fu_1970_p2);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage14 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_pp0_stage15 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_pp0_stage16 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_pp0_stage17 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_pp0_stage18 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_pp0_stage19 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage20 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_pp0_stage21 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_pp0_stage22 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_pp0_stage23 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_pp0_stage24 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_pp0_stage25 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_pp0_stage26 = ap_CS_fsm[32'd26];

    assign ap_CS_fsm_pp0_stage27 = ap_CS_fsm[32'd27];

    assign ap_CS_fsm_pp0_stage28 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_pp0_stage29 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage30 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_pp0_stage31 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_pp0_stage32 = ap_CS_fsm[32'd32];

    assign ap_CS_fsm_pp0_stage33 = ap_CS_fsm[32'd33];

    assign ap_CS_fsm_pp0_stage34 = ap_CS_fsm[32'd34];

    assign ap_CS_fsm_pp0_stage35 = ap_CS_fsm[32'd35];

    assign ap_CS_fsm_pp0_stage36 = ap_CS_fsm[32'd36];

    assign ap_CS_fsm_pp0_stage38 = ap_CS_fsm[32'd38];

    assign ap_CS_fsm_pp0_stage39 = ap_CS_fsm[32'd39];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage40 = ap_CS_fsm[32'd40];

    assign ap_CS_fsm_pp0_stage41 = ap_CS_fsm[32'd41];

    assign ap_CS_fsm_pp0_stage42 = ap_CS_fsm[32'd42];

    assign ap_CS_fsm_pp0_stage43 = ap_CS_fsm[32'd43];

    assign ap_CS_fsm_pp0_stage44 = ap_CS_fsm[32'd44];

    assign ap_CS_fsm_pp0_stage45 = ap_CS_fsm[32'd45];

    assign ap_CS_fsm_pp0_stage46 = ap_CS_fsm[32'd46];

    assign ap_CS_fsm_pp0_stage47 = ap_CS_fsm[32'd47];

    assign ap_CS_fsm_pp0_stage48 = ap_CS_fsm[32'd48];

    assign ap_CS_fsm_pp0_stage49 = ap_CS_fsm[32'd49];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage50 = ap_CS_fsm[32'd50];

    assign ap_CS_fsm_pp0_stage51 = ap_CS_fsm[32'd51];

    assign ap_CS_fsm_pp0_stage52 = ap_CS_fsm[32'd52];

    assign ap_CS_fsm_pp0_stage53 = ap_CS_fsm[32'd53];

    assign ap_CS_fsm_pp0_stage54 = ap_CS_fsm[32'd54];

    assign ap_CS_fsm_pp0_stage55 = ap_CS_fsm[32'd55];

    assign ap_CS_fsm_pp0_stage56 = ap_CS_fsm[32'd56];

    assign ap_CS_fsm_pp0_stage57 = ap_CS_fsm[32'd57];

    assign ap_CS_fsm_pp0_stage58 = ap_CS_fsm[32'd58];

    assign ap_CS_fsm_pp0_stage59 = ap_CS_fsm[32'd59];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage60 = ap_CS_fsm[32'd60];

    assign ap_CS_fsm_pp0_stage61 = ap_CS_fsm[32'd61];

    assign ap_CS_fsm_pp0_stage62 = ap_CS_fsm[32'd62];

    assign ap_CS_fsm_pp0_stage63 = ap_CS_fsm[32'd63];

    assign ap_CS_fsm_pp0_stage64 = ap_CS_fsm[32'd64];

    assign ap_CS_fsm_pp0_stage65 = ap_CS_fsm[32'd65];

    assign ap_CS_fsm_pp0_stage66 = ap_CS_fsm[32'd66];

    assign ap_CS_fsm_pp0_stage67 = ap_CS_fsm[32'd67];

    assign ap_CS_fsm_pp0_stage68 = ap_CS_fsm[32'd68];

    assign ap_CS_fsm_pp0_stage69 = ap_CS_fsm[32'd69];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage70 = ap_CS_fsm[32'd70];

    assign ap_CS_fsm_pp0_stage71 = ap_CS_fsm[32'd71];

    assign ap_CS_fsm_pp0_stage72 = ap_CS_fsm[32'd72];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage53 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage53_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage53_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage54 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage54_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage54_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage55 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage55_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage55_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage56 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage56_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage56_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage57 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage57_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage57_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage58 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage58_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage58_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage59 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage59_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage59_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage60 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage60_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage60_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage61 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage61_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage61_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage62 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage62_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage62_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage63 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage63_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage64 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage64_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage65 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage65_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage66_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage66_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage67 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage67_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage67_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage68 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage68_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage68_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage69 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage69_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage69_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage70_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage70_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage71_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage71_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage72_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    always @(*) begin
        ap_condition_2356 = ((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22));
    end

    always @(*) begin
        ap_condition_3574 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58));
    end

    always @(*) begin
        ap_condition_3579 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage58) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage58));
    end

    always @(*) begin
        ap_condition_3586 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46));
    end

    always @(*) begin
        ap_condition_3591 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage46) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage46));
    end

    always @(*) begin
        ap_condition_3597 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59));
    end

    always @(*) begin
        ap_condition_3602 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage59) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage59));
    end

    always @(*) begin
        ap_condition_3607 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24));
    end

    always @(*) begin
        ap_condition_3612 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage24) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage24));
    end

    always @(*) begin
        ap_condition_3618 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage52) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage52));
    end

    always @(*) begin
        ap_condition_3623 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage52) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage52));
    end

    always @(*) begin
        ap_condition_3629 = ((icmp_ln263_reg_3394 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53));
    end

    always @(*) begin
        ap_condition_3634 = ((icmp_ln263_reg_3394 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage53) & (icmp_ln218_reg_3292 == 1'd0) & (1'b0 == ap_block_pp0_stage53));
    end

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage23;

    always @(*) begin
        ap_predicate_op247_call_state12_state11 = ((1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0));
    end

    always @(*) begin
        ap_predicate_op255_call_state13_state12 = ((1'd1 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0));
    end

    always @(*) begin
        ap_predicate_op321_call_state19_state18 = ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
    end

    always @(*) begin
        ap_predicate_op331_call_state20_state19 = ((((1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_reg_3612) & (1'd1 == and_ln208_5_reg_3697) & (1'd1 == and_ln208_4_reg_3678) & (1'd1 == and_ln208_3_reg_3659) & (icmp_ln218_reg_3292 == 1'd0)));
    end

    always @(*) begin
        ap_predicate_op425_call_state25_state24 = (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
    end

    always @(*) begin
        ap_predicate_op472_call_state26_state25 = (((((((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) & (1'd0 == and_ln208_2_reg_3650) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_5_reg_3697) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_4_reg_3678) & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0))) | ((1'd0 == and_ln208_3_reg_3659) 
    & (1'd0 == and_ln208_1_reg_3631) & (1'd1 == and_ln208_7_reg_3740) & (1'd1 == and_ln208_6_reg_3721) & (1'd1 == and_ln208_reg_3612) & (icmp_ln218_reg_3292 == 1'd0)));
    end

    assign bitcast_ln208_1_fu_2842_p1 = reg_1977;

    assign bitcast_ln208_2_fu_2882_p1 = reg_1982;

    assign bitcast_ln208_3_fu_2927_p1 = reg_1977;

    assign bitcast_ln208_4_fu_2967_p1 = reg_1982;

    assign bitcast_ln208_5_fu_3007_p1 = reg_1977;

    assign bitcast_ln208_6_fu_3047_p1 = reg_1982;

    assign bitcast_ln208_fu_2801_p1 = l_axis_0_load_reg_3478;

    assign bitcast_ln221_1_fu_3128_p1 = xor_ln221_fu_3122_p2;

    assign bitcast_ln221_fu_3118_p1 = reg_2616;

    assign bitcast_ln237_1_fu_3143_p1 = xor_ln237_fu_3137_p2;

    assign bitcast_ln237_fu_3133_p1 = reg_2616;

    assign bitcast_ln251_1_fu_3158_p1 = xor_ln251_fu_3152_p2;

    assign bitcast_ln251_fu_3148_p1 = reg_2616;

    assign grp_sin_or_cos_double_s_fu_1842_ap_start = grp_sin_or_cos_double_s_fu_1842_ap_start_reg;

    assign icmp_ln208_10_fu_3025_p2 = ((tmp_282_fu_3011_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_11_fu_3031_p2 = ((trunc_ln208_5_fu_3021_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_12_fu_3065_p2 = ((tmp_284_fu_3051_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_13_fu_3071_p2 = ((trunc_ln208_6_fu_3061_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_1_fu_2824_p2 = ((trunc_ln208_fu_2814_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_2_fu_2860_p2 = ((tmp_273_fu_2846_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_3_fu_2866_p2 = ((trunc_ln208_1_fu_2856_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_4_fu_2900_p2 = ((tmp_275_fu_2886_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_5_fu_2906_p2 = ((trunc_ln208_2_fu_2896_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_6_fu_2945_p2 = ((tmp_278_fu_2931_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_7_fu_2951_p2 = ((trunc_ln208_3_fu_2941_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_8_fu_2985_p2 = ((tmp_280_fu_2971_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln208_9_fu_2991_p2 = ((trunc_ln208_4_fu_2981_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln208_fu_2818_p2 = ((tmp_271_fu_2804_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln218_fu_2768_p2 = ((ap_sig_allocacmp_idx_5 == 3'd6) ? 1'b1 : 1'b0);

    assign icmp_ln263_fu_2795_p2 = ((ap_sig_allocacmp_idx_5 == 3'd0) ? 1'b1 : 1'b0);

    assign l_axis_0_address0 = zext_ln218_fu_2774_p1;

    assign l_axis_1_addr_1_gep_fu_562_p3 = zext_ln218_reg_3296;

    assign l_axis_1_addr_2_gep_fu_746_p3 = zext_ln218_reg_3296;

    assign l_axis_2_addr_1_gep_fu_738_p3 = zext_ln218_reg_3296;

    assign l_axis_2_addr_2_gep_fu_876_p3 = zext_ln218_reg_3296;

    assign or_ln208_1_fu_2872_p2 = (icmp_ln208_3_reg_3626 | icmp_ln208_2_reg_3621);

    assign or_ln208_2_fu_2912_p2 = (icmp_ln208_5_reg_3645 | icmp_ln208_4_reg_3640);

    assign or_ln208_3_fu_2957_p2 = (icmp_ln208_7_reg_3673 | icmp_ln208_6_reg_3668);

    assign or_ln208_4_fu_2997_p2 = (icmp_ln208_9_reg_3692 | icmp_ln208_8_reg_3687);

    assign or_ln208_5_fu_3037_p2 = (icmp_ln208_11_reg_3716 | icmp_ln208_10_reg_3711);

    assign or_ln208_6_fu_3077_p2 = (icmp_ln208_13_reg_3735 | icmp_ln208_12_reg_3730);

    assign or_ln208_fu_2830_p2 = (icmp_ln208_fu_2818_p2 | icmp_ln208_1_fu_2824_p2);

    assign this_TCurr_0_0_d0 = reg_2451;

    assign this_TCurr_0_2_d0 = reg_2451;

    assign this_TCurr_1_2_d0 = reg_2462;

    assign this_TCurr_2_2_d0 = reg_2475;

    assign this_TCurr_3_2_d0 = reg_2488;

    assign this_TJoint_0_0_addr_1_gep_fu_1321_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_0_addr_3_gep_fu_1470_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_0_addr_4_gep_fu_1518_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_1_addr_1_gep_fu_1337_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_1_addr_3_gep_fu_892_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_1_addr_4_gep_fu_1377_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_2_addr_2_gep_fu_790_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_2_addr_3_gep_fu_1502_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_2_addr_4_gep_fu_1560_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_3_addr_2_gep_fu_798_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_3_addr_3_gep_fu_900_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_3_addr_4_gep_fu_1282_p3 = zext_ln218_reg_3296;

    assign this_TJoint_0_3_d0 = 64'd0;

    assign this_TJoint_1_0_addr_1_gep_fu_1345_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_0_addr_3_gep_fu_908_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_0_addr_4_gep_fu_1369_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_1_addr_1_gep_fu_1329_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_1_addr_2_gep_fu_1387_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_1_addr_4_gep_fu_1427_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_2_addr_2_gep_fu_1411_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_2_addr_3_gep_fu_930_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_2_addr_4_gep_fu_1460_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_3_addr_2_gep_fu_820_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_3_addr_3_gep_fu_938_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_3_addr_4_gep_fu_1290_p3 = zext_ln218_reg_3296;

    assign this_TJoint_1_3_d0 = 64'd0;

    assign this_TJoint_2_0_addr_2_gep_fu_828_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_0_addr_3_gep_fu_1510_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_0_addr_4_gep_fu_1552_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_1_addr_2_gep_fu_1419_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_1_addr_3_gep_fu_946_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_1_addr_4_gep_fu_1452_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_2_addr_2_gep_fu_1395_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_2_addr_3_gep_fu_1478_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_2_addr_4_gep_fu_1526_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_3_addr_2_gep_fu_836_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_3_addr_3_gep_fu_954_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_3_addr_4_gep_fu_1298_p3 = zext_ln218_reg_3296;

    assign this_TJoint_2_3_d0 = 64'd0;

    assign this_TJoint_3_0_addr_2_gep_fu_844_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_0_addr_3_gep_fu_962_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_0_addr_4_gep_fu_1258_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_0_d0 = 64'd0;

    assign this_TJoint_3_1_addr_2_gep_fu_852_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_1_addr_3_gep_fu_970_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_1_addr_4_gep_fu_1266_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_1_d0 = 64'd0;

    assign this_TJoint_3_2_addr_2_gep_fu_860_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_2_addr_3_gep_fu_978_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_2_addr_4_gep_fu_1274_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_2_d0 = 64'd0;

    assign this_TJoint_3_3_addr_2_gep_fu_868_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_3_addr_3_gep_fu_986_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_3_addr_4_gep_fu_1306_p3 = zext_ln218_reg_3296;

    assign this_TJoint_3_3_d0 = 64'd4607182418800017408;

    assign this_TLink_0_0_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_0_1_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_0_2_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_0_3_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_1_0_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_1_1_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_1_2_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_1_3_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_2_0_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_2_1_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_2_2_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_2_3_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_3_0_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_3_1_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_3_2_address0 = zext_ln218_fu_2774_p1;

    assign this_TLink_3_3_address0 = zext_ln218_fu_2774_p1;

    assign this_q_addr_1_gep_fu_754_p3 = zext_ln218_reg_3296;

    assign this_q_addr_2_gep_fu_884_p3 = zext_ln218_reg_3296;

    assign tmp_271_fu_2804_p4 = {{bitcast_ln208_fu_2801_p1[62:52]}};

    assign tmp_273_fu_2846_p4 = {{bitcast_ln208_1_fu_2842_p1[62:52]}};

    assign tmp_275_fu_2886_p4 = {{bitcast_ln208_2_fu_2882_p1[62:52]}};

    assign tmp_278_fu_2931_p4 = {{bitcast_ln208_3_fu_2927_p1[62:52]}};

    assign tmp_280_fu_2971_p4 = {{bitcast_ln208_4_fu_2967_p1[62:52]}};

    assign tmp_282_fu_3011_p4 = {{bitcast_ln208_5_fu_3007_p1[62:52]}};

    assign tmp_284_fu_3051_p4 = {{bitcast_ln208_6_fu_3047_p1[62:52]}};

    assign trunc_ln208_1_fu_2856_p1 = bitcast_ln208_1_fu_2842_p1[51:0];

    assign trunc_ln208_2_fu_2896_p1 = bitcast_ln208_2_fu_2882_p1[51:0];

    assign trunc_ln208_3_fu_2941_p1 = bitcast_ln208_3_fu_2927_p1[51:0];

    assign trunc_ln208_4_fu_2981_p1 = bitcast_ln208_4_fu_2967_p1[51:0];

    assign trunc_ln208_5_fu_3021_p1 = bitcast_ln208_5_fu_3007_p1[51:0];

    assign trunc_ln208_6_fu_3061_p1 = bitcast_ln208_6_fu_3047_p1[51:0];

    assign trunc_ln208_fu_2814_p1 = bitcast_ln208_fu_2801_p1[51:0];

    assign xor_ln221_fu_3122_p2 = (bitcast_ln221_fu_3118_p1 ^ 64'd9223372036854775808);

    assign xor_ln237_fu_3137_p2 = (bitcast_ln237_fu_3133_p1 ^ 64'd9223372036854775808);

    assign xor_ln251_fu_3152_p2 = (bitcast_ln251_fu_3148_p1 ^ 64'd9223372036854775808);

    assign zext_ln218_fu_2774_p1 = ap_sig_allocacmp_idx_5;

    assign zext_ln37_fu_3097_p1 = add_ln267_fu_3092_p2;

    always @(posedge ap_clk) begin
        zext_ln218_reg_3296[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        zext_ln218_reg_3296_pp0_iter1_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        zext_ln37_reg_3749[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_forwardKin_Pipeline_VITIS_LOOP_218_3
