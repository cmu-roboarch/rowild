/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    invOut_address0,
    invOut_ce0,
    invOut_we0,
    invOut_d0,
    inv_address0,
    inv_ce0,
    inv_q0,
    det
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [3:0] invOut_address0;
    output invOut_ce0;
    output invOut_we0;
    output [63:0] invOut_d0;
    output [3:0] inv_address0;
    output inv_ce0;
    input [63:0] inv_q0;
    input [63:0] det;

    reg ap_idle;
    reg invOut_ce0;
    reg invOut_we0;
    reg inv_ce0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln153_fu_112_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] zext_ln155_1_fu_180_p1;
    reg   [63:0] zext_ln155_1_reg_235;
    wire    ap_block_pp0_stage0;
    reg   [2:0] j_fu_44;
    wire   [2:0] add_ln154_fu_185_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_j_load;
    reg   [2:0] i_fu_48;
    wire   [2:0] select_ln153_1_fu_150_p3;
    reg   [2:0] ap_sig_allocacmp_i_load;
    reg   [4:0] indvar_flatten_fu_52;
    wire   [4:0] add_ln153_1_fu_118_p2;
    reg   [4:0] ap_sig_allocacmp_indvar_flatten_load;
    wire   [63:0] mul_fu_88_p2;
    wire   [0:0] icmp_ln154_fu_136_p2;
    wire   [2:0] add_ln153_fu_130_p2;
    wire   [1:0] trunc_ln155_fu_158_p1;
    wire   [2:0] select_ln153_fu_142_p3;
    wire   [3:0] tmp_4_fu_162_p3;
    wire   [3:0] zext_ln155_fu_170_p1;
    wire   [3:0] add_ln155_fu_174_p2;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 j_fu_44 = 3'd0;
        #0 i_fu_48 = 3'd0;
        #0 indvar_flatten_fu_52 = 5'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U1 (
        .din0(inv_q0),
        .din1(det),
        .dout(mul_fu_88_p2)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln153_fu_112_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                i_fu_48 <= select_ln153_1_fu_150_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                i_fu_48 <= 3'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln153_fu_112_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                indvar_flatten_fu_52 <= add_ln153_1_fu_118_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                indvar_flatten_fu_52 <= 5'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln153_fu_112_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                j_fu_44 <= add_ln154_fu_185_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                j_fu_44 <= 3'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            zext_ln155_1_reg_235[3 : 0] <= zext_ln155_1_fu_180_p1[3 : 0];
        end
    end

    always @(*) begin
        if (((icmp_ln153_fu_112_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_i_load = 3'd0;
        end else begin
            ap_sig_allocacmp_i_load = i_fu_48;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_indvar_flatten_load = 5'd0;
        end else begin
            ap_sig_allocacmp_indvar_flatten_load = indvar_flatten_fu_52;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_j_load = 3'd0;
        end else begin
            ap_sig_allocacmp_j_load = j_fu_44;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            invOut_ce0 = 1'b1;
        end else begin
            invOut_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            invOut_we0 = 1'b1;
        end else begin
            invOut_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            inv_ce0 = 1'b1;
        end else begin
            inv_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln153_1_fu_118_p2 = (ap_sig_allocacmp_indvar_flatten_load + 5'd1);

    assign add_ln153_fu_130_p2 = (ap_sig_allocacmp_i_load + 3'd1);

    assign add_ln154_fu_185_p2 = (select_ln153_fu_142_p3 + 3'd1);

    assign add_ln155_fu_174_p2 = (tmp_4_fu_162_p3 + zext_ln155_fu_170_p1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign icmp_ln153_fu_112_p2 = ((ap_sig_allocacmp_indvar_flatten_load == 5'd16) ? 1'b1 : 1'b0);

    assign icmp_ln154_fu_136_p2 = ((ap_sig_allocacmp_j_load == 3'd4) ? 1'b1 : 1'b0);

    assign invOut_address0 = zext_ln155_1_reg_235;

    assign invOut_d0 = mul_fu_88_p2;

    assign inv_address0 = zext_ln155_1_fu_180_p1;

    assign select_ln153_1_fu_150_p3 = ((icmp_ln154_fu_136_p2[0:0] == 1'b1) ? add_ln153_fu_130_p2 : ap_sig_allocacmp_i_load);

    assign select_ln153_fu_142_p3 = ((icmp_ln154_fu_136_p2[0:0] == 1'b1) ? 3'd0 : ap_sig_allocacmp_j_load);

    assign tmp_4_fu_162_p3 = {{trunc_ln155_fu_158_p1}, {2'd0}};

    assign trunc_ln155_fu_158_p1 = select_ln153_1_fu_150_p3[1:0];

    assign zext_ln155_1_fu_180_p1 = add_ln155_fu_174_p2;

    assign zext_ln155_fu_170_p1 = select_ln153_fu_142_p3;

    always @(posedge ap_clk) begin
        zext_ln155_1_reg_235[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2
