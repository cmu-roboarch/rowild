/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_planRRT_Pipeline_VITIS_LOOP_152_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    lfsr_load,
    qRand_address0,
    qRand_ce0,
    qRand_we0,
    qRand_d0,
    or_i_i_i110_out,
    or_i_i_i110_out_ap_vld,
    shr6_i_i_i_phi_out,
    shr6_i_i_i_phi_out_ap_vld,
    grp_fu_1431_p_din0,
    grp_fu_1431_p_din1,
    grp_fu_1431_p_dout0,
    grp_fu_1431_p_ce,
    grp_fu_1436_p_din0,
    grp_fu_1436_p_dout0,
    grp_fu_1436_p_ce,
    grp_fu_1439_p_din0,
    grp_fu_1439_p_dout0,
    grp_fu_1439_p_ce,
    grp_fu_2529_p_din0,
    grp_fu_2529_p_din1,
    grp_fu_2529_p_opcode,
    grp_fu_2529_p_dout0,
    grp_fu_2529_p_ce,
    grp_fu_2533_p_din0,
    grp_fu_2533_p_din1,
    grp_fu_2533_p_dout0,
    grp_fu_2533_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [15:0] lfsr_load;
    output [2:0] qRand_address0;
    output qRand_ce0;
    output qRand_we0;
    output [63:0] qRand_d0;
    output [15:0] or_i_i_i110_out;
    output or_i_i_i110_out_ap_vld;
    output [5:0] shr6_i_i_i_phi_out;
    output shr6_i_i_i_phi_out_ap_vld;
    output [31:0] grp_fu_1431_p_din0;
    output [31:0] grp_fu_1431_p_din1;
    input [31:0] grp_fu_1431_p_dout0;
    output grp_fu_1431_p_ce;
    output [31:0] grp_fu_1436_p_din0;
    input [31:0] grp_fu_1436_p_dout0;
    output grp_fu_1436_p_ce;
    output [31:0] grp_fu_1439_p_din0;
    input [63:0] grp_fu_1439_p_dout0;
    output grp_fu_1439_p_ce;
    output [63:0] grp_fu_2529_p_din0;
    output [63:0] grp_fu_2529_p_din1;
    output [0:0] grp_fu_2529_p_opcode;
    input [63:0] grp_fu_2529_p_dout0;
    output grp_fu_2529_p_ce;
    output [63:0] grp_fu_2533_p_din0;
    output [63:0] grp_fu_2533_p_din1;
    input [63:0] grp_fu_2533_p_dout0;
    output grp_fu_2533_p_ce;

    reg ap_idle;
    reg qRand_ce0;
    reg qRand_we0;
    reg or_i_i_i110_out_ap_vld;
    reg shr6_i_i_i_phi_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_enable_reg_pp0_iter27;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln152_fu_143_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    reg   [2:0] i_reg_284;
    reg   [2:0] i_reg_284_pp0_iter1_reg;
    reg   [2:0] i_reg_284_pp0_iter2_reg;
    reg   [2:0] i_reg_284_pp0_iter3_reg;
    reg   [2:0] i_reg_284_pp0_iter4_reg;
    reg   [2:0] i_reg_284_pp0_iter5_reg;
    reg   [2:0] i_reg_284_pp0_iter6_reg;
    reg   [2:0] i_reg_284_pp0_iter7_reg;
    reg   [2:0] i_reg_284_pp0_iter8_reg;
    reg   [2:0] i_reg_284_pp0_iter9_reg;
    reg   [2:0] i_reg_284_pp0_iter10_reg;
    reg   [2:0] i_reg_284_pp0_iter11_reg;
    reg   [2:0] i_reg_284_pp0_iter12_reg;
    reg   [2:0] i_reg_284_pp0_iter13_reg;
    reg   [2:0] i_reg_284_pp0_iter14_reg;
    reg   [2:0] i_reg_284_pp0_iter15_reg;
    reg   [2:0] i_reg_284_pp0_iter16_reg;
    reg   [2:0] i_reg_284_pp0_iter17_reg;
    reg   [2:0] i_reg_284_pp0_iter18_reg;
    reg   [2:0] i_reg_284_pp0_iter19_reg;
    reg   [2:0] i_reg_284_pp0_iter20_reg;
    reg   [2:0] i_reg_284_pp0_iter21_reg;
    reg   [2:0] i_reg_284_pp0_iter22_reg;
    reg   [2:0] i_reg_284_pp0_iter23_reg;
    reg   [2:0] i_reg_284_pp0_iter24_reg;
    reg   [2:0] i_reg_284_pp0_iter25_reg;
    reg   [2:0] i_reg_284_pp0_iter26_reg;
    reg   [0:0] icmp_ln152_reg_289;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter1_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter2_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter3_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter4_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter5_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter6_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter7_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter8_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter9_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter10_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter11_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter12_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter13_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter14_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter15_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter16_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter17_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter18_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter19_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter20_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter21_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter22_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter23_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter24_reg;
    reg   [0:0] icmp_ln152_reg_289_pp0_iter25_reg;
    wire   [15:0] rand_int_fu_224_p3;
    reg   [15:0] rand_int_reg_293;
    wire   [31:0] zext_ln47_fu_247_p1;
    reg   [31:0] conv_i_i_reg_303;
    reg   [31:0] div_i_i_reg_308;
    reg   [63:0] r_reg_313;
    reg   [63:0] mul_i_reg_318;
    reg   [63:0] add_i_reg_323;
    wire   [63:0] zext_ln152_fu_251_p1;
    wire    ap_block_pp0_stage0;
    reg   [5:0] shr6_i_i_i_phi_fu_64;
    reg   [2:0] i_1_fu_68;
    wire   [2:0] add_ln152_fu_149_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_i;
    reg   [15:0] or_i_i_i110_fu_72;
    reg   [15:0] ap_sig_allocacmp_or_i_i_i110_load;
    wire    ap_block_pp0_stage0_01001;
    wire   [0:0] tmp_14_fu_170_p3;
    wire   [0:0] tmp_15_fu_178_p3;
    wire   [0:0] xor_ln38_fu_206_p2;
    wire   [0:0] tmp_fu_162_p3;
    wire   [0:0] xor_ln38_2_fu_212_p2;
    wire   [0:0] trunc_ln37_fu_158_p1;
    wire   [0:0] xor_ln38_1_fu_218_p2;
    wire   [14:0] lshr_ln38_1_fu_186_p4;
    wire    ap_block_pp0_stage0_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg    ap_loop_exit_ready_pp0_iter10_reg;
    reg    ap_loop_exit_ready_pp0_iter11_reg;
    reg    ap_loop_exit_ready_pp0_iter12_reg;
    reg    ap_loop_exit_ready_pp0_iter13_reg;
    reg    ap_loop_exit_ready_pp0_iter14_reg;
    reg    ap_loop_exit_ready_pp0_iter15_reg;
    reg    ap_loop_exit_ready_pp0_iter16_reg;
    reg    ap_loop_exit_ready_pp0_iter17_reg;
    reg    ap_loop_exit_ready_pp0_iter18_reg;
    reg    ap_loop_exit_ready_pp0_iter19_reg;
    reg    ap_loop_exit_ready_pp0_iter20_reg;
    reg    ap_loop_exit_ready_pp0_iter21_reg;
    reg    ap_loop_exit_ready_pp0_iter22_reg;
    reg    ap_loop_exit_ready_pp0_iter23_reg;
    reg    ap_loop_exit_ready_pp0_iter24_reg;
    reg    ap_loop_exit_ready_pp0_iter25_reg;
    reg    ap_loop_exit_ready_pp0_iter26_reg;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter27 = 1'b0;
        #0 shr6_i_i_i_phi_fu_64 = 6'd0;
        #0 i_1_fu_68 = 3'd0;
        #0 or_i_i_i110_fu_72 = 16'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready_pp0_iter26_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter27 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln152_fu_143_p2 == 1'd0))) begin
                i_1_fu_68 <= add_ln152_fu_149_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                i_1_fu_68 <= 3'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln152_fu_143_p2 == 1'd0))) begin
                or_i_i_i110_fu_72 <= rand_int_fu_224_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                or_i_i_i110_fu_72 <= lfsr_load;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            add_i_reg_323 <= grp_fu_2529_p_dout0;
            ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
            ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
            ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
            ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
            ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
            ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
            ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
            ap_loop_exit_ready_pp0_iter17_reg <= ap_loop_exit_ready_pp0_iter16_reg;
            ap_loop_exit_ready_pp0_iter18_reg <= ap_loop_exit_ready_pp0_iter17_reg;
            ap_loop_exit_ready_pp0_iter19_reg <= ap_loop_exit_ready_pp0_iter18_reg;
            ap_loop_exit_ready_pp0_iter20_reg <= ap_loop_exit_ready_pp0_iter19_reg;
            ap_loop_exit_ready_pp0_iter21_reg <= ap_loop_exit_ready_pp0_iter20_reg;
            ap_loop_exit_ready_pp0_iter22_reg <= ap_loop_exit_ready_pp0_iter21_reg;
            ap_loop_exit_ready_pp0_iter23_reg <= ap_loop_exit_ready_pp0_iter22_reg;
            ap_loop_exit_ready_pp0_iter24_reg <= ap_loop_exit_ready_pp0_iter23_reg;
            ap_loop_exit_ready_pp0_iter25_reg <= ap_loop_exit_ready_pp0_iter24_reg;
            ap_loop_exit_ready_pp0_iter26_reg <= ap_loop_exit_ready_pp0_iter25_reg;
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
            conv_i_i_reg_303 <= grp_fu_1436_p_dout0;
            div_i_i_reg_308 <= grp_fu_1431_p_dout0;
            i_reg_284_pp0_iter10_reg <= i_reg_284_pp0_iter9_reg;
            i_reg_284_pp0_iter11_reg <= i_reg_284_pp0_iter10_reg;
            i_reg_284_pp0_iter12_reg <= i_reg_284_pp0_iter11_reg;
            i_reg_284_pp0_iter13_reg <= i_reg_284_pp0_iter12_reg;
            i_reg_284_pp0_iter14_reg <= i_reg_284_pp0_iter13_reg;
            i_reg_284_pp0_iter15_reg <= i_reg_284_pp0_iter14_reg;
            i_reg_284_pp0_iter16_reg <= i_reg_284_pp0_iter15_reg;
            i_reg_284_pp0_iter17_reg <= i_reg_284_pp0_iter16_reg;
            i_reg_284_pp0_iter18_reg <= i_reg_284_pp0_iter17_reg;
            i_reg_284_pp0_iter19_reg <= i_reg_284_pp0_iter18_reg;
            i_reg_284_pp0_iter20_reg <= i_reg_284_pp0_iter19_reg;
            i_reg_284_pp0_iter21_reg <= i_reg_284_pp0_iter20_reg;
            i_reg_284_pp0_iter22_reg <= i_reg_284_pp0_iter21_reg;
            i_reg_284_pp0_iter23_reg <= i_reg_284_pp0_iter22_reg;
            i_reg_284_pp0_iter24_reg <= i_reg_284_pp0_iter23_reg;
            i_reg_284_pp0_iter25_reg <= i_reg_284_pp0_iter24_reg;
            i_reg_284_pp0_iter26_reg <= i_reg_284_pp0_iter25_reg;
            i_reg_284_pp0_iter2_reg <= i_reg_284_pp0_iter1_reg;
            i_reg_284_pp0_iter3_reg <= i_reg_284_pp0_iter2_reg;
            i_reg_284_pp0_iter4_reg <= i_reg_284_pp0_iter3_reg;
            i_reg_284_pp0_iter5_reg <= i_reg_284_pp0_iter4_reg;
            i_reg_284_pp0_iter6_reg <= i_reg_284_pp0_iter5_reg;
            i_reg_284_pp0_iter7_reg <= i_reg_284_pp0_iter6_reg;
            i_reg_284_pp0_iter8_reg <= i_reg_284_pp0_iter7_reg;
            i_reg_284_pp0_iter9_reg <= i_reg_284_pp0_iter8_reg;
            icmp_ln152_reg_289_pp0_iter10_reg <= icmp_ln152_reg_289_pp0_iter9_reg;
            icmp_ln152_reg_289_pp0_iter11_reg <= icmp_ln152_reg_289_pp0_iter10_reg;
            icmp_ln152_reg_289_pp0_iter12_reg <= icmp_ln152_reg_289_pp0_iter11_reg;
            icmp_ln152_reg_289_pp0_iter13_reg <= icmp_ln152_reg_289_pp0_iter12_reg;
            icmp_ln152_reg_289_pp0_iter14_reg <= icmp_ln152_reg_289_pp0_iter13_reg;
            icmp_ln152_reg_289_pp0_iter15_reg <= icmp_ln152_reg_289_pp0_iter14_reg;
            icmp_ln152_reg_289_pp0_iter16_reg <= icmp_ln152_reg_289_pp0_iter15_reg;
            icmp_ln152_reg_289_pp0_iter17_reg <= icmp_ln152_reg_289_pp0_iter16_reg;
            icmp_ln152_reg_289_pp0_iter18_reg <= icmp_ln152_reg_289_pp0_iter17_reg;
            icmp_ln152_reg_289_pp0_iter19_reg <= icmp_ln152_reg_289_pp0_iter18_reg;
            icmp_ln152_reg_289_pp0_iter20_reg <= icmp_ln152_reg_289_pp0_iter19_reg;
            icmp_ln152_reg_289_pp0_iter21_reg <= icmp_ln152_reg_289_pp0_iter20_reg;
            icmp_ln152_reg_289_pp0_iter22_reg <= icmp_ln152_reg_289_pp0_iter21_reg;
            icmp_ln152_reg_289_pp0_iter23_reg <= icmp_ln152_reg_289_pp0_iter22_reg;
            icmp_ln152_reg_289_pp0_iter24_reg <= icmp_ln152_reg_289_pp0_iter23_reg;
            icmp_ln152_reg_289_pp0_iter25_reg <= icmp_ln152_reg_289_pp0_iter24_reg;
            icmp_ln152_reg_289_pp0_iter2_reg <= icmp_ln152_reg_289_pp0_iter1_reg;
            icmp_ln152_reg_289_pp0_iter3_reg <= icmp_ln152_reg_289_pp0_iter2_reg;
            icmp_ln152_reg_289_pp0_iter4_reg <= icmp_ln152_reg_289_pp0_iter3_reg;
            icmp_ln152_reg_289_pp0_iter5_reg <= icmp_ln152_reg_289_pp0_iter4_reg;
            icmp_ln152_reg_289_pp0_iter6_reg <= icmp_ln152_reg_289_pp0_iter5_reg;
            icmp_ln152_reg_289_pp0_iter7_reg <= icmp_ln152_reg_289_pp0_iter6_reg;
            icmp_ln152_reg_289_pp0_iter8_reg <= icmp_ln152_reg_289_pp0_iter7_reg;
            icmp_ln152_reg_289_pp0_iter9_reg <= icmp_ln152_reg_289_pp0_iter8_reg;
            mul_i_reg_318 <= grp_fu_2533_p_dout0;
            r_reg_313 <= grp_fu_1439_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
            i_reg_284 <= ap_sig_allocacmp_i;
            i_reg_284_pp0_iter1_reg <= i_reg_284;
            icmp_ln152_reg_289 <= icmp_ln152_fu_143_p2;
            icmp_ln152_reg_289_pp0_iter1_reg <= icmp_ln152_reg_289;
            rand_int_reg_293 <= rand_int_fu_224_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln152_fu_143_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            shr6_i_i_i_phi_fu_64 <= {{ap_sig_allocacmp_or_i_i_i110_load[6:1]}};
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln152_fu_143_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready_pp0_iter26_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_idle_pp0 == 1'b1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_i = 3'd0;
        end else begin
            ap_sig_allocacmp_i = i_1_fu_68;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_or_i_i_i110_load = lfsr_load;
        end else begin
            ap_sig_allocacmp_or_i_i_i110_load = or_i_i_i110_fu_72;
        end
    end

    always @(*) begin
        if (((icmp_ln152_reg_289_pp0_iter25_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            or_i_i_i110_out_ap_vld = 1'b1;
        end else begin
            or_i_i_i110_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter27 == 1'b1))) begin
            qRand_ce0 = 1'b1;
        end else begin
            qRand_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter27 == 1'b1))) begin
            qRand_we0 = 1'b1;
        end else begin
            qRand_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln152_reg_289_pp0_iter25_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            shr6_i_i_i_phi_out_ap_vld = 1'b1;
        end else begin
            shr6_i_i_i_phi_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln152_fu_149_p2 = (ap_sig_allocacmp_i + 3'd1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign grp_fu_1431_p_ce = 1'b1;

    assign grp_fu_1431_p_din0 = conv_i_i_reg_303;

    assign grp_fu_1431_p_din1 = 32'd796917760;

    assign grp_fu_1436_p_ce = 1'b1;

    assign grp_fu_1436_p_din0 = zext_ln47_fu_247_p1;

    assign grp_fu_1439_p_ce = 1'b1;

    assign grp_fu_1439_p_din0 = div_i_i_reg_308;

    assign grp_fu_2529_p_ce = 1'b1;

    assign grp_fu_2529_p_din0 = mul_i_reg_318;

    assign grp_fu_2529_p_din1 = 64'd13833125093780374864;

    assign grp_fu_2529_p_opcode = 2'd0;

    assign grp_fu_2533_p_ce = 1'b1;

    assign grp_fu_2533_p_din0 = r_reg_313;

    assign grp_fu_2533_p_din1 = 64'd4614256656552969552;

    assign icmp_ln152_fu_143_p2 = ((ap_sig_allocacmp_i == 3'd5) ? 1'b1 : 1'b0);

    assign lshr_ln38_1_fu_186_p4 = {{ap_sig_allocacmp_or_i_i_i110_load[15:1]}};

    assign or_i_i_i110_out = or_i_i_i110_fu_72;

    assign qRand_address0 = zext_ln152_fu_251_p1;

    assign qRand_d0 = add_i_reg_323;

    assign rand_int_fu_224_p3 = {{xor_ln38_1_fu_218_p2}, {lshr_ln38_1_fu_186_p4}};

    assign shr6_i_i_i_phi_out = shr6_i_i_i_phi_fu_64;

    assign tmp_14_fu_170_p3 = ap_sig_allocacmp_or_i_i_i110_load[32'd2];

    assign tmp_15_fu_178_p3 = ap_sig_allocacmp_or_i_i_i110_load[32'd5];

    assign tmp_fu_162_p3 = ap_sig_allocacmp_or_i_i_i110_load[32'd3];

    assign trunc_ln37_fu_158_p1 = ap_sig_allocacmp_or_i_i_i110_load[0:0];

    assign xor_ln38_1_fu_218_p2 = (xor_ln38_2_fu_212_p2 ^ trunc_ln37_fu_158_p1);

    assign xor_ln38_2_fu_212_p2 = (xor_ln38_fu_206_p2 ^ tmp_fu_162_p3);

    assign xor_ln38_fu_206_p2 = (tmp_15_fu_178_p3 ^ tmp_14_fu_170_p3);

    assign zext_ln152_fu_251_p1 = i_reg_284_pp0_iter26_reg;

    assign zext_ln47_fu_247_p1 = rand_int_reg_293;

endmodule  //main_planRRT_Pipeline_VITIS_LOOP_152_1
