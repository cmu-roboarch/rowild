/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_rayCast (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    pf_address0,
    pf_ce0,
    pf_q0,
    x,
    y,
    theta,
    degree,
    ap_return,
    grp_fu_597_p_din0,
    grp_fu_597_p_din1,
    grp_fu_597_p_opcode,
    grp_fu_597_p_dout0,
    grp_fu_597_p_ce,
    grp_fu_601_p_din0,
    grp_fu_601_p_din1,
    grp_fu_601_p_opcode,
    grp_fu_601_p_dout0,
    grp_fu_601_p_ce,
    grp_fu_605_p_din0,
    grp_fu_605_p_din1,
    grp_fu_605_p_dout0,
    grp_fu_605_p_ce,
    grp_fu_609_p_din0,
    grp_fu_609_p_din1,
    grp_fu_609_p_dout0,
    grp_fu_609_p_ce,
    grp_fu_613_p_din0,
    grp_fu_613_p_dout0,
    grp_fu_613_p_ce,
    grp_fu_616_p_din0,
    grp_fu_616_p_din1,
    grp_fu_616_p_opcode,
    grp_fu_616_p_dout0,
    grp_fu_616_p_ce,
    grp_fu_221_p_din0,
    grp_fu_221_p_din1,
    grp_fu_221_p_dout0,
    grp_fu_221_p_ce,
    grp_fu_620_p_din0,
    grp_fu_620_p_din1,
    grp_fu_620_p_opcode,
    grp_fu_620_p_dout0,
    grp_fu_620_p_ce,
    grp_sin_or_cos_double_s_fu_624_p_din1,
    grp_sin_or_cos_double_s_fu_624_p_din2,
    grp_sin_or_cos_double_s_fu_624_p_dout0,
    grp_sin_or_cos_double_s_fu_624_p_start,
    grp_sin_or_cos_double_s_fu_624_p_ready,
    grp_sin_or_cos_double_s_fu_624_p_done,
    grp_sin_or_cos_double_s_fu_624_p_idle,
    grp_sin_or_cos_double_s_fu_635_p_din1,
    grp_sin_or_cos_double_s_fu_635_p_din2,
    grp_sin_or_cos_double_s_fu_635_p_dout0,
    grp_sin_or_cos_double_s_fu_635_p_start,
    grp_sin_or_cos_double_s_fu_635_p_ready,
    grp_sin_or_cos_double_s_fu_635_p_done,
    grp_sin_or_cos_double_s_fu_635_p_idle
);

    parameter ap_ST_fsm_state1 = 26'd1;
    parameter ap_ST_fsm_state2 = 26'd2;
    parameter ap_ST_fsm_state3 = 26'd4;
    parameter ap_ST_fsm_state4 = 26'd8;
    parameter ap_ST_fsm_state5 = 26'd16;
    parameter ap_ST_fsm_state6 = 26'd32;
    parameter ap_ST_fsm_state7 = 26'd64;
    parameter ap_ST_fsm_state8 = 26'd128;
    parameter ap_ST_fsm_state9 = 26'd256;
    parameter ap_ST_fsm_state10 = 26'd512;
    parameter ap_ST_fsm_state11 = 26'd1024;
    parameter ap_ST_fsm_state12 = 26'd2048;
    parameter ap_ST_fsm_state13 = 26'd4096;
    parameter ap_ST_fsm_state14 = 26'd8192;
    parameter ap_ST_fsm_state15 = 26'd16384;
    parameter ap_ST_fsm_state16 = 26'd32768;
    parameter ap_ST_fsm_state17 = 26'd65536;
    parameter ap_ST_fsm_state18 = 26'd131072;
    parameter ap_ST_fsm_state19 = 26'd262144;
    parameter ap_ST_fsm_state20 = 26'd524288;
    parameter ap_ST_fsm_state21 = 26'd1048576;
    parameter ap_ST_fsm_state22 = 26'd2097152;
    parameter ap_ST_fsm_state23 = 26'd4194304;
    parameter ap_ST_fsm_state24 = 26'd8388608;
    parameter ap_ST_fsm_state25 = 26'd16777216;
    parameter ap_ST_fsm_state26 = 26'd33554432;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [16:0] pf_address0;
    output pf_ce0;
    input [255:0] pf_q0;
    input [63:0] x;
    input [63:0] y;
    input [63:0] theta;
    input [63:0] degree;
    output [63:0] ap_return;
    output [63:0] grp_fu_597_p_din0;
    output [63:0] grp_fu_597_p_din1;
    output [1:0] grp_fu_597_p_opcode;
    input [63:0] grp_fu_597_p_dout0;
    output grp_fu_597_p_ce;
    output [63:0] grp_fu_601_p_din0;
    output [63:0] grp_fu_601_p_din1;
    output [0:0] grp_fu_601_p_opcode;
    input [63:0] grp_fu_601_p_dout0;
    output grp_fu_601_p_ce;
    output [63:0] grp_fu_605_p_din0;
    output [63:0] grp_fu_605_p_din1;
    input [63:0] grp_fu_605_p_dout0;
    output grp_fu_605_p_ce;
    output [63:0] grp_fu_609_p_din0;
    output [63:0] grp_fu_609_p_din1;
    input [63:0] grp_fu_609_p_dout0;
    output grp_fu_609_p_ce;
    output [31:0] grp_fu_613_p_din0;
    input [63:0] grp_fu_613_p_dout0;
    output grp_fu_613_p_ce;
    output [31:0] grp_fu_616_p_din0;
    output [31:0] grp_fu_616_p_din1;
    output [4:0] grp_fu_616_p_opcode;
    input [0:0] grp_fu_616_p_dout0;
    output grp_fu_616_p_ce;
    output [63:0] grp_fu_221_p_din0;
    output [63:0] grp_fu_221_p_din1;
    input [63:0] grp_fu_221_p_dout0;
    output grp_fu_221_p_ce;
    output [63:0] grp_fu_620_p_din0;
    output [63:0] grp_fu_620_p_din1;
    output [4:0] grp_fu_620_p_opcode;
    input [0:0] grp_fu_620_p_dout0;
    output grp_fu_620_p_ce;
    output [63:0] grp_sin_or_cos_double_s_fu_624_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_624_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_624_p_dout0;
    output grp_sin_or_cos_double_s_fu_624_p_start;
    input grp_sin_or_cos_double_s_fu_624_p_ready;
    input grp_sin_or_cos_double_s_fu_624_p_done;
    input grp_sin_or_cos_double_s_fu_624_p_idle;
    output [63:0] grp_sin_or_cos_double_s_fu_635_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_635_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_635_p_dout0;
    output grp_sin_or_cos_double_s_fu_635_p_start;
    input grp_sin_or_cos_double_s_fu_635_p_ready;
    input grp_sin_or_cos_double_s_fu_635_p_done;
    input grp_sin_or_cos_double_s_fu_635_p_idle;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[16:0] pf_address0;
    reg pf_ce0;

    (* fsm_encoding = "none" *) reg   [25:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    reg   [63:0] reg_201;
    wire    ap_CS_fsm_state7;
    wire    ap_CS_fsm_state14;
    wire    ap_CS_fsm_state23;
    reg   [63:0] reg_209;
    wire    ap_CS_fsm_state16;
    reg    ap_block_state16_on_subcall_done;
    reg   [63:0] reg_216;
    wire    ap_CS_fsm_state9;
    reg    ap_block_state9_on_subcall_done;
    reg   [63:0] reg_221;
    reg   [63:0] reg_226;
    wire    ap_CS_fsm_state8;
    reg   [63:0] trunc_ln_reg_344;
    wire   [63:0] trunc_ln217_fu_242_p1;
    reg   [63:0] trunc_ln217_reg_349;
    wire   [63:0] bitcast_ln214_fu_246_p1;
    wire    ap_CS_fsm_state10;
    wire    ap_CS_fsm_state17;
    wire   [63:0] step_fu_251_p1;
    reg   [63:0] step_reg_370;
    wire    ap_CS_fsm_state22;
    reg   [63:0] yRay_reg_382;
    wire   [190:0] empty_fu_256_p1;
    reg   [190:0] empty_reg_387;
    reg   [63:0] p_cast_reg_392;
    reg   [63:0] trunc_ln3_reg_397;
    reg   [10:0] tmp_30_reg_402;
    reg   [51:0] trunc_ln230_1_reg_407;
    reg   [51:0] trunc_ln235_3_reg_412;
    wire   [63:0] empty_70_fu_310_p1;
    reg   [63:0] empty_70_reg_417;
    wire    ap_CS_fsm_state24;
    wire   [63:0] bitcast_ln235_fu_314_p1;
    reg   [63:0] bitcast_ln235_reg_422;
    wire    grp_sin_or_cos_double_s_fu_123_ap_ready;
    reg   [63:0] grp_sin_or_cos_double_s_fu_123_t_in;
    wire    grp_sin_or_cos_double_s_fu_142_ap_ready;
    reg   [63:0] grp_sin_or_cos_double_s_fu_142_t_in;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_done;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_idle;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_ready;
    wire   [16:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_address0;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_ce0;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out_ap_vld;
    wire   [31:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_din0;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_ce;
    wire   [31:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din0;
    wire   [31:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din1;
    wire   [4:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_opcode;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_ce;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din0;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din1;
    wire   [0:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_opcode;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_ce;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din0;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din1;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_ce;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din0;
    wire   [63:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din1;
    wire   [4:0] grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_opcode;
    wire    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_ce;
    reg    grp_sin_or_cos_double_s_fu_123_ap_start_reg;
    wire    ap_CS_fsm_state15;
    reg    grp_sin_or_cos_double_s_fu_142_ap_start_reg;
    reg    grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg;
    wire    ap_CS_fsm_state25;
    reg   [63:0] dist_1_loc_fu_72;
    wire    ap_CS_fsm_state26;
    reg   [63:0] grp_fu_179_p0;
    reg   [63:0] grp_fu_179_p1;
    reg   [63:0] grp_fu_191_p0;
    reg   [63:0] grp_fu_191_p1;
    reg   [63:0] grp_fu_197_p0;
    reg   [1:0] grp_fu_179_opcode;
    reg    grp_fu_179_ce;
    wire    ap_CS_fsm_state2;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    wire    ap_CS_fsm_state5;
    wire    ap_CS_fsm_state6;
    reg    grp_fu_191_ce;
    reg    grp_fu_197_ce;
    reg    grp_fu_427_ce;
    reg    grp_fu_430_ce;
    reg    grp_fu_434_ce;
    reg    grp_fu_438_ce;
    reg   [25:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    reg    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    reg    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    reg    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 26'd1;
        #0 grp_sin_or_cos_double_s_fu_123_ap_start_reg = 1'b0;
        #0 grp_sin_or_cos_double_s_fu_142_ap_start_reg = 1'b0;
        #0 grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg = 1'b0;
    end

    main_rayCast_Pipeline_VITIS_LOOP_222_1 grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start),
        .ap_done(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_done),
        .ap_idle(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_idle),
        .ap_ready(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_ready),
        .xRay(reg_201),
        .yRay(yRay_reg_382),
        .step(step_reg_370),
        .xStep(reg_209),
        .yStep(reg_226),
        .tmp_30(tmp_30_reg_402),
        .trunc_ln230_1(trunc_ln230_1_reg_407),
        .empty(empty_70_reg_417),
        .pf_address0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_address0),
        .pf_ce0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_ce0),
        .pf_q0(pf_q0),
        .pf_load_6(empty_reg_387),
        .trunc_ln235_3(trunc_ln235_3_reg_412),
        .bitcast_ln235(bitcast_ln235_reg_422),
        .dist_1_out(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out),
        .dist_1_out_ap_vld(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out_ap_vld),
        .grp_fu_427_p_din0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_din0),
        .grp_fu_427_p_dout0(grp_fu_613_p_dout0),
        .grp_fu_427_p_ce(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_ce),
        .grp_fu_430_p_din0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din0),
        .grp_fu_430_p_din1(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din1),
        .grp_fu_430_p_opcode(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_opcode),
        .grp_fu_430_p_dout0(grp_fu_616_p_dout0),
        .grp_fu_430_p_ce(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_ce),
        .grp_fu_179_p_din0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din0),
        .grp_fu_179_p_din1(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din1),
        .grp_fu_179_p_opcode(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_opcode),
        .grp_fu_179_p_dout0(grp_fu_597_p_dout0),
        .grp_fu_179_p_ce(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_ce),
        .grp_fu_434_p_din0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din0),
        .grp_fu_434_p_din1(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din1),
        .grp_fu_434_p_dout0(grp_fu_221_p_dout0),
        .grp_fu_434_p_ce(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_ce),
        .grp_fu_438_p_din0(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din0),
        .grp_fu_438_p_din1(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din1),
        .grp_fu_438_p_opcode(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_opcode),
        .grp_fu_438_p_dout0(grp_fu_620_p_dout0),
        .grp_fu_438_p_ce(grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_ce)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state24)) begin
                grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg <= 1'b1;
            end else if ((grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_ready == 1'b1)) begin
                grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_123_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state8))) begin
                grp_sin_or_cos_double_s_fu_123_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_123_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_123_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_142_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state8))) begin
                grp_sin_or_cos_double_s_fu_142_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_142_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_142_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state24)) begin
            bitcast_ln235_reg_422 <= bitcast_ln235_fu_314_p1;
            empty_70_reg_417 <= empty_70_fu_310_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state25))) begin
            dist_1_loc_fu_72 <= grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_dist_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state23)) begin
            empty_reg_387 <= empty_fu_256_p1;
            p_cast_reg_392 <= {{pf_q0[255:192]}};
            tmp_30_reg_402 <= {{pf_q0[254:244]}};
            trunc_ln230_1_reg_407 <= {{pf_q0[243:192]}};
            trunc_ln235_3_reg_412 <= {{pf_q0[179:128]}};
            trunc_ln3_reg_397 <= {{pf_q0[191:128]}};
            yRay_reg_382 <= grp_fu_601_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state7))) begin
            reg_201 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state7) | ((1'b0 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16)))) begin
            reg_209 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16)) | ((1'b0 == ap_block_state9_on_subcall_done) & (1'b1 == ap_CS_fsm_state9)))) begin
            reg_216 <= grp_sin_or_cos_double_s_fu_624_p_dout0;
            reg_221 <= grp_sin_or_cos_double_s_fu_635_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state23) | ((1'b0 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16)))) begin
            reg_226 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            step_reg_370 <= step_fu_251_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            trunc_ln217_reg_349 <= trunc_ln217_fu_242_p1;
            trunc_ln_reg_344 <= {{pf_q0[127:64]}};
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state16_on_subcall_done)) begin
            ap_ST_fsm_state16_blk = 1'b1;
        end else begin
            ap_ST_fsm_state16_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    always @(*) begin
        if ((grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_done == 1'b0)) begin
            ap_ST_fsm_state25_blk = 1'b1;
        end else begin
            ap_ST_fsm_state25_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state9_on_subcall_done)) begin
            ap_ST_fsm_state9_blk = 1'b1;
        end else begin
            ap_ST_fsm_state9_blk = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state26) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state26)) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_179_ce = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_ce;
        end else if (((1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state24) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) | ((1'b1 == ap_block_state9_on_subcall_done) & (1'b1 == ap_CS_fsm_state9)))) begin
            grp_fu_179_ce = 1'b0;
        end else begin
            grp_fu_179_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_179_opcode = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_179_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state17) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
            grp_fu_179_opcode = 2'd0;
        end else begin
            grp_fu_179_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_179_p0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_179_p0 = reg_209;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_179_p0 = reg_201;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_179_p0 = theta;
        end else begin
            grp_fu_179_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_179_p1 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_179_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_179_p1 = x;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_179_p1 = reg_209;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_179_p1 = 64'd4609753056925599056;
        end else begin
            grp_fu_179_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9) | ((1'b1 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16)) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            grp_fu_191_ce = 1'b0;
        end else begin
            grp_fu_191_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_191_p0 = step_fu_251_p1;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_191_p0 = bitcast_ln214_fu_246_p1;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_191_p0 = degree;
        end else begin
            grp_fu_191_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state10))) begin
            grp_fu_191_p1 = reg_216;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_191_p1 = 64'd4580687790477189905;
        end else begin
            grp_fu_191_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state1) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9) | ((1'b1 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16)))) begin
            grp_fu_197_ce = 1'b0;
        end else begin
            grp_fu_197_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_197_p0 = step_fu_251_p1;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_197_p0 = bitcast_ln214_fu_246_p1;
        end else begin
            grp_fu_197_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_427_ce = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_ce;
        end else begin
            grp_fu_427_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_430_ce = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_ce;
        end else begin
            grp_fu_430_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_434_ce = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_ce;
        end else begin
            grp_fu_434_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state25)) begin
            grp_fu_438_ce = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_ce;
        end else begin
            grp_fu_438_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state16)) begin
            grp_sin_or_cos_double_s_fu_123_t_in = reg_201;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_sin_or_cos_double_s_fu_123_t_in = theta;
        end else begin
            grp_sin_or_cos_double_s_fu_123_t_in = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state16)) begin
            grp_sin_or_cos_double_s_fu_142_t_in = reg_201;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_sin_or_cos_double_s_fu_142_t_in = theta;
        end else begin
            grp_sin_or_cos_double_s_fu_142_t_in = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state22)) begin
            pf_address0 = 64'd80502;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            pf_address0 = 64'd80503;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            pf_address0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_address0;
        end else begin
            pf_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state8))) begin
            pf_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            pf_ce0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_pf_ce0;
        end else begin
            pf_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                if (((1'b0 == ap_block_state9_on_subcall_done) & (1'b1 == ap_CS_fsm_state9))) begin
                    ap_NS_fsm = ap_ST_fsm_state10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state9;
                end
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                if (((1'b0 == ap_block_state16_on_subcall_done) & (1'b1 == ap_CS_fsm_state16))) begin
                    ap_NS_fsm = ap_ST_fsm_state17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state16;
                end
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                if (((1'b1 == ap_CS_fsm_state25) & (grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state26;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state25;
                end
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ap_CS_fsm_state1  = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state2  = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_state3  = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4  = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5  = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6  = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state7  = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state8  = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state9  = ap_CS_fsm[32'd8];

    always @(*) begin
        ap_block_state16_on_subcall_done = ((grp_sin_or_cos_double_s_fu_635_p_done == 1'b0) | (grp_sin_or_cos_double_s_fu_624_p_done == 1'b0));
    end

    always @(*) begin
        ap_block_state9_on_subcall_done = ((grp_sin_or_cos_double_s_fu_635_p_done == 1'b0) | (grp_sin_or_cos_double_s_fu_624_p_done == 1'b0));
    end

    assign ap_return = dist_1_loc_fu_72;

    assign bitcast_ln214_fu_246_p1 = trunc_ln_reg_344;

    assign bitcast_ln235_fu_314_p1 = trunc_ln3_reg_397;

    assign empty_70_fu_310_p1 = p_cast_reg_392;

    assign empty_fu_256_p1 = pf_q0[190:0];

    assign grp_fu_221_p_ce = grp_fu_434_ce;

    assign grp_fu_221_p_din0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din0;

    assign grp_fu_221_p_din1 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_434_p_din1;

    assign grp_fu_597_p_ce = grp_fu_179_ce;

    assign grp_fu_597_p_din0 = grp_fu_179_p0;

    assign grp_fu_597_p_din1 = grp_fu_179_p1;

    assign grp_fu_597_p_opcode = grp_fu_179_opcode;

    assign grp_fu_601_p_ce = 1'b1;

    assign grp_fu_601_p_din0 = reg_226;

    assign grp_fu_601_p_din1 = y;

    assign grp_fu_601_p_opcode = 2'd0;

    assign grp_fu_605_p_ce = grp_fu_191_ce;

    assign grp_fu_605_p_din0 = grp_fu_191_p0;

    assign grp_fu_605_p_din1 = grp_fu_191_p1;

    assign grp_fu_609_p_ce = grp_fu_197_ce;

    assign grp_fu_609_p_din0 = grp_fu_197_p0;

    assign grp_fu_609_p_din1 = reg_221;

    assign grp_fu_613_p_ce = grp_fu_427_ce;

    assign grp_fu_613_p_din0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_427_p_din0;

    assign grp_fu_616_p_ce = grp_fu_430_ce;

    assign grp_fu_616_p_din0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din0;

    assign grp_fu_616_p_din1 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_din1;

    assign grp_fu_616_p_opcode = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_430_p_opcode;

    assign grp_fu_620_p_ce = grp_fu_438_ce;

    assign grp_fu_620_p_din0 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din0;

    assign grp_fu_620_p_din1 = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_din1;

    assign grp_fu_620_p_opcode = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_grp_fu_438_p_opcode;

    assign grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start = grp_rayCast_Pipeline_VITIS_LOOP_222_1_fu_161_ap_start_reg;

    assign grp_sin_or_cos_double_s_fu_123_ap_ready = grp_sin_or_cos_double_s_fu_624_p_ready;

    assign grp_sin_or_cos_double_s_fu_142_ap_ready = grp_sin_or_cos_double_s_fu_635_p_ready;

    assign grp_sin_or_cos_double_s_fu_624_p_din1 = grp_sin_or_cos_double_s_fu_123_t_in;

    assign grp_sin_or_cos_double_s_fu_624_p_din2 = 1'd1;

    assign grp_sin_or_cos_double_s_fu_624_p_start = grp_sin_or_cos_double_s_fu_123_ap_start_reg;

    assign grp_sin_or_cos_double_s_fu_635_p_din1 = grp_sin_or_cos_double_s_fu_142_t_in;

    assign grp_sin_or_cos_double_s_fu_635_p_din2 = 1'd0;

    assign grp_sin_or_cos_double_s_fu_635_p_start = grp_sin_or_cos_double_s_fu_142_ap_start_reg;

    assign step_fu_251_p1 = trunc_ln217_reg_349;

    assign trunc_ln217_fu_242_p1 = pf_q0[63:0];

endmodule  //main_rayCast
