/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_38_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    env_axesObs_address0,
    env_axesObs_ce0,
    env_axesObs_we0,
    env_axesObs_d0,
    env_axesObs_address1,
    env_axesObs_ce1,
    env_axesObs_we1,
    env_axesObs_d1,
    env_pointsObs_0_0_address0,
    env_pointsObs_0_0_ce0,
    env_pointsObs_0_0_we0,
    env_pointsObs_0_0_d0,
    env_pointsObs_0_1_address0,
    env_pointsObs_0_1_ce0,
    env_pointsObs_0_1_we0,
    env_pointsObs_0_1_d0,
    env_pointsObs_0_2_address0,
    env_pointsObs_0_2_ce0,
    env_pointsObs_0_2_we0,
    env_pointsObs_0_2_d0,
    env_pointsObs_1_0_address0,
    env_pointsObs_1_0_ce0,
    env_pointsObs_1_0_we0,
    env_pointsObs_1_0_d0,
    env_pointsObs_1_1_address0,
    env_pointsObs_1_1_ce0,
    env_pointsObs_1_1_we0,
    env_pointsObs_1_1_d0,
    env_pointsObs_1_2_address0,
    env_pointsObs_1_2_ce0,
    env_pointsObs_1_2_we0,
    env_pointsObs_1_2_d0,
    env_pointsObs_2_0_address0,
    env_pointsObs_2_0_ce0,
    env_pointsObs_2_0_we0,
    env_pointsObs_2_0_d0,
    env_pointsObs_2_1_address0,
    env_pointsObs_2_1_ce0,
    env_pointsObs_2_1_we0,
    env_pointsObs_2_1_d0,
    env_pointsObs_2_2_address0,
    env_pointsObs_2_2_ce0,
    env_pointsObs_2_2_we0,
    env_pointsObs_2_2_d0,
    env_pointsObs_3_0_address0,
    env_pointsObs_3_0_ce0,
    env_pointsObs_3_0_we0,
    env_pointsObs_3_0_d0,
    env_pointsObs_3_1_address0,
    env_pointsObs_3_1_ce0,
    env_pointsObs_3_1_we0,
    env_pointsObs_3_1_d0,
    env_pointsObs_3_2_address0,
    env_pointsObs_3_2_ce0,
    env_pointsObs_3_2_we0,
    env_pointsObs_3_2_d0,
    env_pointsObs_4_0_address0,
    env_pointsObs_4_0_ce0,
    env_pointsObs_4_0_we0,
    env_pointsObs_4_0_d0,
    env_pointsObs_4_1_address0,
    env_pointsObs_4_1_ce0,
    env_pointsObs_4_1_we0,
    env_pointsObs_4_1_d0,
    env_pointsObs_4_2_address0,
    env_pointsObs_4_2_ce0,
    env_pointsObs_4_2_we0,
    env_pointsObs_4_2_d0,
    env_pointsObs_5_0_address0,
    env_pointsObs_5_0_ce0,
    env_pointsObs_5_0_we0,
    env_pointsObs_5_0_d0,
    env_pointsObs_5_1_address0,
    env_pointsObs_5_1_ce0,
    env_pointsObs_5_1_we0,
    env_pointsObs_5_1_d0,
    env_pointsObs_5_2_address0,
    env_pointsObs_5_2_ce0,
    env_pointsObs_5_2_we0,
    env_pointsObs_5_2_d0,
    env_pointsObs_6_0_address0,
    env_pointsObs_6_0_ce0,
    env_pointsObs_6_0_we0,
    env_pointsObs_6_0_d0,
    env_pointsObs_6_1_address0,
    env_pointsObs_6_1_ce0,
    env_pointsObs_6_1_we0,
    env_pointsObs_6_1_d0,
    env_pointsObs_6_2_address0,
    env_pointsObs_6_2_ce0,
    env_pointsObs_6_2_we0,
    env_pointsObs_6_2_d0,
    env_pointsObs_7_0_address0,
    env_pointsObs_7_0_ce0,
    env_pointsObs_7_0_we0,
    env_pointsObs_7_0_d0,
    env_pointsObs_7_1_address0,
    env_pointsObs_7_1_ce0,
    env_pointsObs_7_1_we0,
    env_pointsObs_7_1_d0,
    env_pointsObs_7_2_address0,
    env_pointsObs_7_2_ce0,
    env_pointsObs_7_2_we0,
    env_pointsObs_7_2_d0,
    env_pointsObs_8_0_address0,
    env_pointsObs_8_0_ce0,
    env_pointsObs_8_0_we0,
    env_pointsObs_8_0_d0,
    env_pointsObs_8_1_address0,
    env_pointsObs_8_1_ce0,
    env_pointsObs_8_1_we0,
    env_pointsObs_8_1_d0,
    env_pointsObs_8_2_address0,
    env_pointsObs_8_2_ce0,
    env_pointsObs_8_2_we0,
    env_pointsObs_8_2_d0,
    grp_fu_2403_p_din0,
    grp_fu_2403_p_din1,
    grp_fu_2403_p_opcode,
    grp_fu_2403_p_dout0,
    grp_fu_2403_p_ce,
    grp_fu_2407_p_din0,
    grp_fu_2407_p_din1,
    grp_fu_2407_p_opcode,
    grp_fu_2407_p_dout0,
    grp_fu_2407_p_ce,
    grp_fu_2411_p_din0,
    grp_fu_2411_p_din1,
    grp_fu_2411_p_opcode,
    grp_fu_2411_p_dout0,
    grp_fu_2411_p_ce,
    grp_fu_2415_p_din0,
    grp_fu_2415_p_din1,
    grp_fu_2415_p_opcode,
    grp_fu_2415_p_dout0,
    grp_fu_2415_p_ce,
    grp_fu_2419_p_din0,
    grp_fu_2419_p_din1,
    grp_fu_2419_p_opcode,
    grp_fu_2419_p_dout0,
    grp_fu_2419_p_ce,
    grp_fu_2423_p_din0,
    grp_fu_2423_p_din1,
    grp_fu_2423_p_opcode,
    grp_fu_2423_p_dout0,
    grp_fu_2423_p_ce,
    grp_fu_2427_p_din0,
    grp_fu_2427_p_din1,
    grp_fu_2427_p_opcode,
    grp_fu_2427_p_dout0,
    grp_fu_2427_p_ce,
    grp_fu_2431_p_din0,
    grp_fu_2431_p_din1,
    grp_fu_2431_p_dout0,
    grp_fu_2431_p_ce,
    grp_fu_2435_p_din0,
    grp_fu_2435_p_din1,
    grp_fu_2435_p_dout0,
    grp_fu_2435_p_ce,
    grp_fu_2439_p_din0,
    grp_fu_2439_p_din1,
    grp_fu_2439_p_dout0,
    grp_fu_2439_p_ce,
    grp_fu_2443_p_din0,
    grp_fu_2443_p_din1,
    grp_fu_2443_p_dout0,
    grp_fu_2443_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 5'd1;
    parameter ap_ST_fsm_pp0_stage1 = 5'd2;
    parameter ap_ST_fsm_pp0_stage2 = 5'd4;
    parameter ap_ST_fsm_pp0_stage3 = 5'd8;
    parameter ap_ST_fsm_pp0_stage4 = 5'd16;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] env_axesObs_address0;
    output env_axesObs_ce0;
    output env_axesObs_we0;
    output [63:0] env_axesObs_d0;
    output [6:0] env_axesObs_address1;
    output env_axesObs_ce1;
    output env_axesObs_we1;
    output [63:0] env_axesObs_d1;
    output [2:0] env_pointsObs_0_0_address0;
    output env_pointsObs_0_0_ce0;
    output env_pointsObs_0_0_we0;
    output [63:0] env_pointsObs_0_0_d0;
    output [2:0] env_pointsObs_0_1_address0;
    output env_pointsObs_0_1_ce0;
    output env_pointsObs_0_1_we0;
    output [63:0] env_pointsObs_0_1_d0;
    output [2:0] env_pointsObs_0_2_address0;
    output env_pointsObs_0_2_ce0;
    output env_pointsObs_0_2_we0;
    output [63:0] env_pointsObs_0_2_d0;
    output [2:0] env_pointsObs_1_0_address0;
    output env_pointsObs_1_0_ce0;
    output env_pointsObs_1_0_we0;
    output [63:0] env_pointsObs_1_0_d0;
    output [2:0] env_pointsObs_1_1_address0;
    output env_pointsObs_1_1_ce0;
    output env_pointsObs_1_1_we0;
    output [63:0] env_pointsObs_1_1_d0;
    output [2:0] env_pointsObs_1_2_address0;
    output env_pointsObs_1_2_ce0;
    output env_pointsObs_1_2_we0;
    output [63:0] env_pointsObs_1_2_d0;
    output [2:0] env_pointsObs_2_0_address0;
    output env_pointsObs_2_0_ce0;
    output env_pointsObs_2_0_we0;
    output [63:0] env_pointsObs_2_0_d0;
    output [2:0] env_pointsObs_2_1_address0;
    output env_pointsObs_2_1_ce0;
    output env_pointsObs_2_1_we0;
    output [63:0] env_pointsObs_2_1_d0;
    output [2:0] env_pointsObs_2_2_address0;
    output env_pointsObs_2_2_ce0;
    output env_pointsObs_2_2_we0;
    output [63:0] env_pointsObs_2_2_d0;
    output [2:0] env_pointsObs_3_0_address0;
    output env_pointsObs_3_0_ce0;
    output env_pointsObs_3_0_we0;
    output [63:0] env_pointsObs_3_0_d0;
    output [2:0] env_pointsObs_3_1_address0;
    output env_pointsObs_3_1_ce0;
    output env_pointsObs_3_1_we0;
    output [63:0] env_pointsObs_3_1_d0;
    output [2:0] env_pointsObs_3_2_address0;
    output env_pointsObs_3_2_ce0;
    output env_pointsObs_3_2_we0;
    output [63:0] env_pointsObs_3_2_d0;
    output [2:0] env_pointsObs_4_0_address0;
    output env_pointsObs_4_0_ce0;
    output env_pointsObs_4_0_we0;
    output [63:0] env_pointsObs_4_0_d0;
    output [2:0] env_pointsObs_4_1_address0;
    output env_pointsObs_4_1_ce0;
    output env_pointsObs_4_1_we0;
    output [63:0] env_pointsObs_4_1_d0;
    output [2:0] env_pointsObs_4_2_address0;
    output env_pointsObs_4_2_ce0;
    output env_pointsObs_4_2_we0;
    output [63:0] env_pointsObs_4_2_d0;
    output [2:0] env_pointsObs_5_0_address0;
    output env_pointsObs_5_0_ce0;
    output env_pointsObs_5_0_we0;
    output [63:0] env_pointsObs_5_0_d0;
    output [2:0] env_pointsObs_5_1_address0;
    output env_pointsObs_5_1_ce0;
    output env_pointsObs_5_1_we0;
    output [63:0] env_pointsObs_5_1_d0;
    output [2:0] env_pointsObs_5_2_address0;
    output env_pointsObs_5_2_ce0;
    output env_pointsObs_5_2_we0;
    output [63:0] env_pointsObs_5_2_d0;
    output [2:0] env_pointsObs_6_0_address0;
    output env_pointsObs_6_0_ce0;
    output env_pointsObs_6_0_we0;
    output [63:0] env_pointsObs_6_0_d0;
    output [2:0] env_pointsObs_6_1_address0;
    output env_pointsObs_6_1_ce0;
    output env_pointsObs_6_1_we0;
    output [63:0] env_pointsObs_6_1_d0;
    output [2:0] env_pointsObs_6_2_address0;
    output env_pointsObs_6_2_ce0;
    output env_pointsObs_6_2_we0;
    output [63:0] env_pointsObs_6_2_d0;
    output [2:0] env_pointsObs_7_0_address0;
    output env_pointsObs_7_0_ce0;
    output env_pointsObs_7_0_we0;
    output [63:0] env_pointsObs_7_0_d0;
    output [2:0] env_pointsObs_7_1_address0;
    output env_pointsObs_7_1_ce0;
    output env_pointsObs_7_1_we0;
    output [63:0] env_pointsObs_7_1_d0;
    output [2:0] env_pointsObs_7_2_address0;
    output env_pointsObs_7_2_ce0;
    output env_pointsObs_7_2_we0;
    output [63:0] env_pointsObs_7_2_d0;
    output [2:0] env_pointsObs_8_0_address0;
    output env_pointsObs_8_0_ce0;
    output env_pointsObs_8_0_we0;
    output [63:0] env_pointsObs_8_0_d0;
    output [2:0] env_pointsObs_8_1_address0;
    output env_pointsObs_8_1_ce0;
    output env_pointsObs_8_1_we0;
    output [63:0] env_pointsObs_8_1_d0;
    output [2:0] env_pointsObs_8_2_address0;
    output env_pointsObs_8_2_ce0;
    output env_pointsObs_8_2_we0;
    output [63:0] env_pointsObs_8_2_d0;
    output [63:0] grp_fu_2403_p_din0;
    output [63:0] grp_fu_2403_p_din1;
    output [1:0] grp_fu_2403_p_opcode;
    input [63:0] grp_fu_2403_p_dout0;
    output grp_fu_2403_p_ce;
    output [63:0] grp_fu_2407_p_din0;
    output [63:0] grp_fu_2407_p_din1;
    output [1:0] grp_fu_2407_p_opcode;
    input [63:0] grp_fu_2407_p_dout0;
    output grp_fu_2407_p_ce;
    output [63:0] grp_fu_2411_p_din0;
    output [63:0] grp_fu_2411_p_din1;
    output [1:0] grp_fu_2411_p_opcode;
    input [63:0] grp_fu_2411_p_dout0;
    output grp_fu_2411_p_ce;
    output [63:0] grp_fu_2415_p_din0;
    output [63:0] grp_fu_2415_p_din1;
    output [1:0] grp_fu_2415_p_opcode;
    input [63:0] grp_fu_2415_p_dout0;
    output grp_fu_2415_p_ce;
    output [63:0] grp_fu_2419_p_din0;
    output [63:0] grp_fu_2419_p_din1;
    output [1:0] grp_fu_2419_p_opcode;
    input [63:0] grp_fu_2419_p_dout0;
    output grp_fu_2419_p_ce;
    output [63:0] grp_fu_2423_p_din0;
    output [63:0] grp_fu_2423_p_din1;
    output [1:0] grp_fu_2423_p_opcode;
    input [63:0] grp_fu_2423_p_dout0;
    output grp_fu_2423_p_ce;
    output [63:0] grp_fu_2427_p_din0;
    output [63:0] grp_fu_2427_p_din1;
    output [1:0] grp_fu_2427_p_opcode;
    input [63:0] grp_fu_2427_p_dout0;
    output grp_fu_2427_p_ce;
    output [63:0] grp_fu_2431_p_din0;
    output [63:0] grp_fu_2431_p_din1;
    input [63:0] grp_fu_2431_p_dout0;
    output grp_fu_2431_p_ce;
    output [63:0] grp_fu_2435_p_din0;
    output [63:0] grp_fu_2435_p_din1;
    input [63:0] grp_fu_2435_p_dout0;
    output grp_fu_2435_p_ce;
    output [63:0] grp_fu_2439_p_din0;
    output [63:0] grp_fu_2439_p_din1;
    input [63:0] grp_fu_2439_p_dout0;
    output grp_fu_2439_p_ce;
    output [63:0] grp_fu_2443_p_din0;
    output [63:0] grp_fu_2443_p_din1;
    input [63:0] grp_fu_2443_p_dout0;
    output grp_fu_2443_p_ce;

    reg ap_idle;
    reg[6:0] env_axesObs_address0;
    reg env_axesObs_ce0;
    reg env_axesObs_we0;
    reg[63:0] env_axesObs_d0;
    reg[6:0] env_axesObs_address1;
    reg env_axesObs_ce1;
    reg env_axesObs_we1;
    reg[63:0] env_axesObs_d1;
    reg env_pointsObs_0_0_ce0;
    reg env_pointsObs_0_0_we0;
    reg env_pointsObs_0_1_ce0;
    reg env_pointsObs_0_1_we0;
    reg env_pointsObs_0_2_ce0;
    reg env_pointsObs_0_2_we0;
    reg env_pointsObs_1_0_ce0;
    reg env_pointsObs_1_0_we0;
    reg env_pointsObs_1_1_ce0;
    reg env_pointsObs_1_1_we0;
    reg env_pointsObs_1_2_ce0;
    reg env_pointsObs_1_2_we0;
    reg env_pointsObs_2_0_ce0;
    reg env_pointsObs_2_0_we0;
    reg env_pointsObs_2_1_ce0;
    reg env_pointsObs_2_1_we0;
    reg env_pointsObs_2_2_ce0;
    reg env_pointsObs_2_2_we0;
    reg env_pointsObs_3_0_ce0;
    reg env_pointsObs_3_0_we0;
    reg env_pointsObs_3_1_ce0;
    reg env_pointsObs_3_1_we0;
    reg env_pointsObs_3_2_ce0;
    reg env_pointsObs_3_2_we0;
    reg env_pointsObs_4_0_ce0;
    reg env_pointsObs_4_0_we0;
    reg env_pointsObs_4_1_ce0;
    reg env_pointsObs_4_1_we0;
    reg env_pointsObs_4_2_ce0;
    reg env_pointsObs_4_2_we0;
    reg env_pointsObs_5_0_ce0;
    reg env_pointsObs_5_0_we0;
    reg env_pointsObs_5_1_ce0;
    reg env_pointsObs_5_1_we0;
    reg env_pointsObs_5_2_ce0;
    reg env_pointsObs_5_2_we0;
    reg env_pointsObs_6_0_ce0;
    reg env_pointsObs_6_0_we0;
    reg env_pointsObs_6_1_ce0;
    reg env_pointsObs_6_1_we0;
    reg env_pointsObs_6_2_ce0;
    reg env_pointsObs_6_2_we0;
    reg env_pointsObs_7_0_ce0;
    reg env_pointsObs_7_0_we0;
    reg env_pointsObs_7_1_ce0;
    reg env_pointsObs_7_1_we0;
    reg env_pointsObs_7_2_ce0;
    reg env_pointsObs_7_2_we0;
    reg env_pointsObs_8_0_ce0;
    reg env_pointsObs_8_0_we0;
    reg env_pointsObs_8_1_ce0;
    reg env_pointsObs_8_1_we0;
    reg env_pointsObs_8_2_ce0;
    reg env_pointsObs_8_2_we0;

    (* fsm_encoding = "none" *) reg   [4:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_subdone;
    reg   [0:0] icmp_ln38_reg_867;
    reg    ap_condition_exit_pp0_iter0_stage4;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    reg   [63:0] reg_609;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    reg   [63:0] reg_615;
    reg   [63:0] reg_621;
    reg   [63:0] reg_627;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] reg_634;
    reg   [63:0] reg_641;
    reg   [63:0] reg_648;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire   [63:0] grp_fu_577_p2;
    reg   [63:0] reg_655;
    wire   [63:0] grp_fu_581_p2;
    reg   [63:0] reg_662;
    reg   [3:0] o_1_reg_860;
    reg   [3:0] o_1_reg_860_pp0_iter1_reg;
    reg   [3:0] o_1_reg_860_pp0_iter2_reg;
    reg   [3:0] o_1_reg_860_pp0_iter3_reg;
    reg   [3:0] o_1_reg_860_pp0_iter4_reg;
    reg   [3:0] o_1_reg_860_pp0_iter5_reg;
    reg   [3:0] o_1_reg_860_pp0_iter6_reg;
    reg   [3:0] o_1_reg_860_pp0_iter7_reg;
    reg   [3:0] o_1_reg_860_pp0_iter8_reg;
    reg   [3:0] o_1_reg_860_pp0_iter9_reg;
    reg   [3:0] o_1_reg_860_pp0_iter10_reg;
    reg   [3:0] o_1_reg_860_pp0_iter11_reg;
    reg   [3:0] o_1_reg_860_pp0_iter12_reg;
    reg   [3:0] o_1_reg_860_pp0_iter13_reg;
    reg   [3:0] o_1_reg_860_pp0_iter14_reg;
    reg   [3:0] o_1_reg_860_pp0_iter15_reg;
    reg   [3:0] o_1_reg_860_pp0_iter16_reg;
    reg   [3:0] o_1_reg_860_pp0_iter17_reg;
    reg   [3:0] o_1_reg_860_pp0_iter18_reg;
    wire   [0:0] icmp_ln38_fu_677_p2;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter1_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter2_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter3_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter4_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter5_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter6_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter7_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter8_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter9_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter10_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter11_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter12_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter13_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter14_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter15_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter16_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter17_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter18_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter19_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter20_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter21_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter22_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter23_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter24_reg;
    reg   [0:0] icmp_ln38_reg_867_pp0_iter25_reg;
    wire   [3:0] indvars_iv_next29_i_fu_683_p2;
    reg   [3:0] indvars_iv_next29_i_reg_871;
    wire   [63:0] grp_fu_606_p1;
    reg   [63:0] conv_i_reg_882;
    reg   [63:0] nums_6_reg_887;
    reg   [63:0] nums_6_reg_887_pp0_iter3_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter4_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter5_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter6_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter7_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter8_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter9_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter10_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter11_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter12_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter13_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter14_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter15_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter16_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter17_reg;
    reg   [63:0] nums_6_reg_887_pp0_iter18_reg;
    reg   [63:0] H_0_0_reg_896;
    reg   [63:0] H_0_1_reg_902;
    reg   [63:0] H_0_2_reg_908;
    reg   [63:0] H_0_3_reg_914;
    reg   [63:0] H_0_3_reg_914_pp0_iter19_reg;
    reg   [63:0] H_0_3_reg_914_pp0_iter20_reg;
    reg   [63:0] H_1_0_reg_921;
    reg   [63:0] H_1_1_reg_927;
    reg   [63:0] H_1_2_reg_933;
    reg   [63:0] H_1_3_reg_939;
    reg   [63:0] H_1_3_reg_939_pp0_iter19_reg;
    reg   [63:0] H_1_3_reg_939_pp0_iter20_reg;
    reg   [63:0] H_2_0_reg_946;
    reg   [63:0] H_2_1_reg_952;
    reg   [63:0] H_2_2_reg_958;
    reg   [63:0] H_2_3_reg_964;
    reg   [63:0] H_2_3_reg_964_pp0_iter19_reg;
    reg   [63:0] H_2_3_reg_964_pp0_iter20_reg;
    wire   [63:0] zext_ln38_fu_745_p1;
    reg   [63:0] zext_ln38_reg_971;
    reg   [63:0] zext_ln38_reg_971_pp0_iter19_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter20_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter21_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter22_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter23_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter24_reg;
    reg   [63:0] zext_ln38_reg_971_pp0_iter25_reg;
    wire   [6:0] add_ln64_fu_761_p2;
    reg   [6:0] add_ln64_reg_999;
    reg   [63:0] mul_i_reg_1010;
    reg   [63:0] mul6_i_reg_1015;
    reg   [63:0] mul3_i_reg_1020;
    reg   [63:0] mul4_i_reg_1025;
    wire    ap_block_pp0_stage4_11001;
    reg   [63:0] mul5_i_reg_1030;
    reg   [63:0] mul7_i_reg_1035;
    reg   [63:0] mul8_i_reg_1040;
    reg   [63:0] mul9_i_reg_1045;
    reg   [63:0] mul1_i_reg_1050;
    reg   [63:0] xL_reg_1055;
    reg   [63:0] xL_1_reg_1061;
    reg   [63:0] xL_2_reg_1067;
    reg   [63:0] yL_reg_1073;
    reg   [63:0] yL_reg_1073_pp0_iter22_reg;
    reg   [63:0] yL_1_reg_1080;
    reg   [63:0] yL_1_reg_1080_pp0_iter22_reg;
    reg   [63:0] yL_2_reg_1087;
    reg   [63:0] yL_2_reg_1087_pp0_iter22_reg;
    reg   [63:0] zL_reg_1094;
    reg   [63:0] zL_reg_1094_pp0_iter22_reg;
    reg   [63:0] zL_reg_1094_pp0_iter23_reg;
    reg   [63:0] zL_reg_1094_pp0_iter24_reg;
    reg   [63:0] zL_1_reg_1101;
    reg   [63:0] zL_1_reg_1101_pp0_iter22_reg;
    reg   [63:0] zL_1_reg_1101_pp0_iter23_reg;
    reg   [63:0] zL_1_reg_1101_pp0_iter24_reg;
    reg   [63:0] zL_2_reg_1108;
    reg   [63:0] zL_2_reg_1108_pp0_iter23_reg;
    reg   [63:0] zL_2_reg_1108_pp0_iter24_reg;
    reg   [63:0] add_i_reg_1115;
    reg   [63:0] add_1_i_reg_1121;
    reg   [63:0] add_2_i_reg_1127;
    reg   [63:0] sub5_i_reg_1133;
    reg   [63:0] sub155_1_i_reg_1139;
    reg   [63:0] sub155_2_i_reg_1145;
    reg   [63:0] add2_i_reg_1151;
    reg   [63:0] add67_1_i_reg_1157;
    reg   [63:0] add67_2_i_reg_1163;
    reg   [63:0] sub3_i_reg_1169;
    reg   [63:0] sub112_1_i_reg_1174;
    reg   [63:0] sub112_2_i_reg_1179;
    reg   [63:0] add5_i_reg_1184;
    reg   [63:0] add158_1_i_reg_1190;
    reg   [63:0] add158_2_i_reg_1196;
    reg   [63:0] sub7_i_reg_1202;
    reg   [63:0] sub204_1_i_reg_1208;
    reg   [63:0] sub204_2_i_reg_1214;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage1_subdone;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_0;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_1;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_2;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_3;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_4;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_5;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_6;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_7;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_8;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_9;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_10;
    wire   [63:0] grp_rpyxyzToH_double_2_fu_544_ap_return_11;
    wire    ap_block_pp0_stage4;
    wire   [63:0] zext_ln64_1_fu_767_p1;
    wire    ap_block_pp0_stage2;
    wire   [63:0] zext_ln64_2_fu_778_p1;
    wire   [63:0] zext_ln64_3_fu_788_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln64_4_fu_798_p1;
    wire   [63:0] zext_ln64_5_fu_808_p1;
    wire   [63:0] zext_ln64_6_fu_818_p1;
    wire   [63:0] zext_ln64_7_fu_828_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln64_8_fu_838_p1;
    wire   [63:0] zext_ln64_9_fu_848_p1;
    wire    ap_block_pp0_stage1;
    reg   [3:0] o_fu_108;
    wire    ap_loop_init;
    reg   [3:0] ap_sig_allocacmp_o_1;
    reg   [63:0] grp_fu_549_p0;
    reg   [63:0] grp_fu_549_p1;
    reg   [63:0] grp_fu_553_p0;
    reg   [63:0] grp_fu_553_p1;
    reg   [63:0] grp_fu_557_p0;
    reg   [63:0] grp_fu_557_p1;
    reg   [63:0] grp_fu_561_p0;
    reg   [63:0] grp_fu_561_p1;
    reg   [63:0] grp_fu_565_p0;
    reg   [63:0] grp_fu_565_p1;
    reg   [63:0] grp_fu_569_p0;
    reg   [63:0] grp_fu_569_p1;
    reg   [63:0] grp_fu_573_p0;
    reg   [63:0] grp_fu_573_p1;
    reg   [63:0] grp_fu_577_p0;
    reg   [63:0] grp_fu_577_p1;
    reg   [63:0] grp_fu_581_p0;
    reg   [63:0] grp_fu_581_p1;
    reg   [63:0] grp_fu_585_p0;
    reg   [63:0] grp_fu_585_p1;
    reg   [63:0] grp_fu_590_p0;
    reg   [63:0] grp_fu_590_p1;
    reg   [63:0] grp_fu_594_p0;
    reg   [63:0] grp_fu_594_p1;
    reg   [63:0] grp_fu_598_p0;
    reg   [63:0] grp_fu_598_p1;
    wire   [31:0] grp_fu_606_p0;
    wire   [6:0] tmp_37_fu_754_p3;
    wire   [6:0] zext_ln64_fu_751_p1;
    wire   [6:0] add_ln64_1_fu_772_p2;
    wire   [6:0] add_ln64_2_fu_783_p2;
    wire   [6:0] add_ln64_3_fu_793_p2;
    wire   [6:0] add_ln64_4_fu_803_p2;
    wire   [6:0] add_ln64_5_fu_813_p2;
    wire   [6:0] add_ln64_6_fu_823_p2;
    wire   [6:0] add_ln64_7_fu_833_p2;
    wire   [6:0] add_ln64_8_fu_843_p2;
    reg   [1:0] grp_fu_549_opcode;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage4_00001;
    reg   [1:0] grp_fu_553_opcode;
    reg   [1:0] grp_fu_557_opcode;
    reg   [1:0] grp_fu_573_opcode;
    reg   [1:0] grp_fu_577_opcode;
    reg   [1:0] grp_fu_581_opcode;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_condition_exit_pp0_iter25_stage1;
    reg    ap_idle_pp0_0to24;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg    ap_loop_exit_ready_pp0_iter10_reg;
    reg    ap_loop_exit_ready_pp0_iter11_reg;
    reg    ap_loop_exit_ready_pp0_iter12_reg;
    reg    ap_loop_exit_ready_pp0_iter13_reg;
    reg    ap_loop_exit_ready_pp0_iter14_reg;
    reg    ap_loop_exit_ready_pp0_iter15_reg;
    reg    ap_loop_exit_ready_pp0_iter16_reg;
    reg    ap_loop_exit_ready_pp0_iter17_reg;
    reg    ap_loop_exit_ready_pp0_iter18_reg;
    reg    ap_loop_exit_ready_pp0_iter19_reg;
    reg    ap_loop_exit_ready_pp0_iter20_reg;
    reg    ap_loop_exit_ready_pp0_iter21_reg;
    reg    ap_loop_exit_ready_pp0_iter22_reg;
    reg    ap_loop_exit_ready_pp0_iter23_reg;
    reg    ap_loop_exit_ready_pp0_iter24_reg;
    reg    ap_loop_exit_ready_pp0_iter25_reg;
    reg   [4:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to26;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 5'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 o_fu_108 = 4'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_rpyxyzToH_double_2 grp_rpyxyzToH_double_2_fu_544 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .x(nums_6_reg_887),
        .ap_return_0(grp_rpyxyzToH_double_2_fu_544_ap_return_0),
        .ap_return_1(grp_rpyxyzToH_double_2_fu_544_ap_return_1),
        .ap_return_2(grp_rpyxyzToH_double_2_fu_544_ap_return_2),
        .ap_return_3(grp_rpyxyzToH_double_2_fu_544_ap_return_3),
        .ap_return_4(grp_rpyxyzToH_double_2_fu_544_ap_return_4),
        .ap_return_5(grp_rpyxyzToH_double_2_fu_544_ap_return_5),
        .ap_return_6(grp_rpyxyzToH_double_2_fu_544_ap_return_6),
        .ap_return_7(grp_rpyxyzToH_double_2_fu_544_ap_return_7),
        .ap_return_8(grp_rpyxyzToH_double_2_fu_544_ap_return_8),
        .ap_return_9(grp_rpyxyzToH_double_2_fu_544_ap_return_9),
        .ap_return_10(grp_rpyxyzToH_double_2_fu_544_ap_return_10),
        .ap_return_11(grp_rpyxyzToH_double_2_fu_544_ap_return_11)
    );

    main_dadddsub_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_U113 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_577_p0),
        .din1(grp_fu_577_p1),
        .opcode(grp_fu_577_opcode),
        .ce(1'b1),
        .dout(grp_fu_577_p2)
    );

    main_dadddsub_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_U114 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_581_p0),
        .din1(grp_fu_581_p1),
        .opcode(grp_fu_581_opcode),
        .ce(1'b1),
        .dout(grp_fu_581_p2)
    );

    main_sitodp_32ns_64_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) sitodp_32ns_64_6_no_dsp_1_U119 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_606_p0),
        .ce(1'b1),
        .dout(grp_fu_606_p1)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage4),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_loop_exit_ready_pp0_iter25_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage4)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
                ap_enable_reg_pp0_iter26 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter17_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter17_reg <= ap_loop_exit_ready_pp0_iter16_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter18_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter18_reg <= ap_loop_exit_ready_pp0_iter17_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter19_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter19_reg <= ap_loop_exit_ready_pp0_iter18_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter20_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter20_reg <= ap_loop_exit_ready_pp0_iter19_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter21_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter21_reg <= ap_loop_exit_ready_pp0_iter20_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter22_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter22_reg <= ap_loop_exit_ready_pp0_iter21_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter23_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter23_reg <= ap_loop_exit_ready_pp0_iter22_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter24_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter24_reg <= ap_loop_exit_ready_pp0_iter23_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter25_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter25_reg <= ap_loop_exit_ready_pp0_iter24_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            o_fu_108 <= 4'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln38_reg_867 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            o_fu_108 <= indvars_iv_next29_i_reg_871;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            H_0_0_reg_896 <= grp_rpyxyzToH_double_2_fu_544_ap_return_0;
            H_0_1_reg_902 <= grp_rpyxyzToH_double_2_fu_544_ap_return_1;
            H_0_2_reg_908 <= grp_rpyxyzToH_double_2_fu_544_ap_return_2;
            H_0_3_reg_914 <= grp_rpyxyzToH_double_2_fu_544_ap_return_3;
            H_0_3_reg_914_pp0_iter19_reg <= H_0_3_reg_914;
            H_0_3_reg_914_pp0_iter20_reg <= H_0_3_reg_914_pp0_iter19_reg;
            H_1_0_reg_921 <= grp_rpyxyzToH_double_2_fu_544_ap_return_4;
            H_1_1_reg_927 <= grp_rpyxyzToH_double_2_fu_544_ap_return_5;
            H_1_2_reg_933 <= grp_rpyxyzToH_double_2_fu_544_ap_return_6;
            H_1_3_reg_939 <= grp_rpyxyzToH_double_2_fu_544_ap_return_7;
            H_1_3_reg_939_pp0_iter19_reg <= H_1_3_reg_939;
            H_1_3_reg_939_pp0_iter20_reg <= H_1_3_reg_939_pp0_iter19_reg;
            H_2_0_reg_946 <= grp_rpyxyzToH_double_2_fu_544_ap_return_8;
            H_2_1_reg_952 <= grp_rpyxyzToH_double_2_fu_544_ap_return_9;
            H_2_2_reg_958 <= grp_rpyxyzToH_double_2_fu_544_ap_return_10;
            H_2_3_reg_964 <= grp_rpyxyzToH_double_2_fu_544_ap_return_11;
            H_2_3_reg_964_pp0_iter19_reg <= H_2_3_reg_964;
            H_2_3_reg_964_pp0_iter20_reg <= H_2_3_reg_964_pp0_iter19_reg;
            conv_i_reg_882 <= grp_fu_606_p1;
            yL_1_reg_1080_pp0_iter22_reg <= yL_1_reg_1080;
            yL_2_reg_1087_pp0_iter22_reg <= yL_2_reg_1087;
            yL_reg_1073_pp0_iter22_reg <= yL_reg_1073;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter23 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            add158_1_i_reg_1190 <= grp_fu_577_p2;
            add158_2_i_reg_1196 <= grp_fu_581_p2;
            add2_i_reg_1151 <= grp_fu_2403_p_dout0;
            add5_i_reg_1184 <= grp_fu_2427_p_dout0;
            add67_1_i_reg_1157 <= grp_fu_2407_p_dout0;
            add67_2_i_reg_1163 <= grp_fu_2411_p_dout0;
            sub112_1_i_reg_1174 <= grp_fu_2419_p_dout0;
            sub112_2_i_reg_1179 <= grp_fu_2423_p_dout0;
            sub3_i_reg_1169 <= grp_fu_2415_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            add_1_i_reg_1121 <= grp_fu_2407_p_dout0;
            add_2_i_reg_1127 <= grp_fu_2411_p_dout0;
            add_i_reg_1115 <= grp_fu_2403_p_dout0;
            sub155_1_i_reg_1139 <= grp_fu_2419_p_dout0;
            sub155_2_i_reg_1145 <= grp_fu_2423_p_dout0;
            sub5_i_reg_1133 <= grp_fu_2415_p_dout0;
            zL_2_reg_1108 <= grp_fu_2439_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            add_ln64_reg_999 <= add_ln64_fu_761_p2;
            zL_1_reg_1101_pp0_iter22_reg <= zL_1_reg_1101;
            zL_1_reg_1101_pp0_iter23_reg <= zL_1_reg_1101_pp0_iter22_reg;
            zL_1_reg_1101_pp0_iter24_reg <= zL_1_reg_1101_pp0_iter23_reg;
            zL_2_reg_1108_pp0_iter23_reg <= zL_2_reg_1108;
            zL_2_reg_1108_pp0_iter24_reg <= zL_2_reg_1108_pp0_iter23_reg;
            zL_reg_1094_pp0_iter22_reg <= zL_reg_1094;
            zL_reg_1094_pp0_iter23_reg <= zL_reg_1094_pp0_iter22_reg;
            zL_reg_1094_pp0_iter24_reg <= zL_reg_1094_pp0_iter23_reg;
            zext_ln38_reg_971[3 : 0] <= zext_ln38_fu_745_p1[3 : 0];
            zext_ln38_reg_971_pp0_iter19_reg[3 : 0] <= zext_ln38_reg_971[3 : 0];
            zext_ln38_reg_971_pp0_iter20_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter19_reg[3 : 0];
            zext_ln38_reg_971_pp0_iter21_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter20_reg[3 : 0];
            zext_ln38_reg_971_pp0_iter22_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter21_reg[3 : 0];
            zext_ln38_reg_971_pp0_iter23_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter22_reg[3 : 0];
            zext_ln38_reg_971_pp0_iter24_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter23_reg[3 : 0];
            zext_ln38_reg_971_pp0_iter25_reg[3 : 0] <= zext_ln38_reg_971_pp0_iter24_reg[3 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            icmp_ln38_reg_867 <= icmp_ln38_fu_677_p2;
            icmp_ln38_reg_867_pp0_iter10_reg <= icmp_ln38_reg_867_pp0_iter9_reg;
            icmp_ln38_reg_867_pp0_iter11_reg <= icmp_ln38_reg_867_pp0_iter10_reg;
            icmp_ln38_reg_867_pp0_iter12_reg <= icmp_ln38_reg_867_pp0_iter11_reg;
            icmp_ln38_reg_867_pp0_iter13_reg <= icmp_ln38_reg_867_pp0_iter12_reg;
            icmp_ln38_reg_867_pp0_iter14_reg <= icmp_ln38_reg_867_pp0_iter13_reg;
            icmp_ln38_reg_867_pp0_iter15_reg <= icmp_ln38_reg_867_pp0_iter14_reg;
            icmp_ln38_reg_867_pp0_iter16_reg <= icmp_ln38_reg_867_pp0_iter15_reg;
            icmp_ln38_reg_867_pp0_iter17_reg <= icmp_ln38_reg_867_pp0_iter16_reg;
            icmp_ln38_reg_867_pp0_iter18_reg <= icmp_ln38_reg_867_pp0_iter17_reg;
            icmp_ln38_reg_867_pp0_iter19_reg <= icmp_ln38_reg_867_pp0_iter18_reg;
            icmp_ln38_reg_867_pp0_iter1_reg <= icmp_ln38_reg_867;
            icmp_ln38_reg_867_pp0_iter20_reg <= icmp_ln38_reg_867_pp0_iter19_reg;
            icmp_ln38_reg_867_pp0_iter21_reg <= icmp_ln38_reg_867_pp0_iter20_reg;
            icmp_ln38_reg_867_pp0_iter22_reg <= icmp_ln38_reg_867_pp0_iter21_reg;
            icmp_ln38_reg_867_pp0_iter23_reg <= icmp_ln38_reg_867_pp0_iter22_reg;
            icmp_ln38_reg_867_pp0_iter24_reg <= icmp_ln38_reg_867_pp0_iter23_reg;
            icmp_ln38_reg_867_pp0_iter25_reg <= icmp_ln38_reg_867_pp0_iter24_reg;
            icmp_ln38_reg_867_pp0_iter2_reg <= icmp_ln38_reg_867_pp0_iter1_reg;
            icmp_ln38_reg_867_pp0_iter3_reg <= icmp_ln38_reg_867_pp0_iter2_reg;
            icmp_ln38_reg_867_pp0_iter4_reg <= icmp_ln38_reg_867_pp0_iter3_reg;
            icmp_ln38_reg_867_pp0_iter5_reg <= icmp_ln38_reg_867_pp0_iter4_reg;
            icmp_ln38_reg_867_pp0_iter6_reg <= icmp_ln38_reg_867_pp0_iter5_reg;
            icmp_ln38_reg_867_pp0_iter7_reg <= icmp_ln38_reg_867_pp0_iter6_reg;
            icmp_ln38_reg_867_pp0_iter8_reg <= icmp_ln38_reg_867_pp0_iter7_reg;
            icmp_ln38_reg_867_pp0_iter9_reg <= icmp_ln38_reg_867_pp0_iter8_reg;
            indvars_iv_next29_i_reg_871 <= indvars_iv_next29_i_fu_683_p2;
            o_1_reg_860 <= ap_sig_allocacmp_o_1;
            o_1_reg_860_pp0_iter10_reg <= o_1_reg_860_pp0_iter9_reg;
            o_1_reg_860_pp0_iter11_reg <= o_1_reg_860_pp0_iter10_reg;
            o_1_reg_860_pp0_iter12_reg <= o_1_reg_860_pp0_iter11_reg;
            o_1_reg_860_pp0_iter13_reg <= o_1_reg_860_pp0_iter12_reg;
            o_1_reg_860_pp0_iter14_reg <= o_1_reg_860_pp0_iter13_reg;
            o_1_reg_860_pp0_iter15_reg <= o_1_reg_860_pp0_iter14_reg;
            o_1_reg_860_pp0_iter16_reg <= o_1_reg_860_pp0_iter15_reg;
            o_1_reg_860_pp0_iter17_reg <= o_1_reg_860_pp0_iter16_reg;
            o_1_reg_860_pp0_iter18_reg <= o_1_reg_860_pp0_iter17_reg;
            o_1_reg_860_pp0_iter1_reg <= o_1_reg_860;
            o_1_reg_860_pp0_iter2_reg <= o_1_reg_860_pp0_iter1_reg;
            o_1_reg_860_pp0_iter3_reg <= o_1_reg_860_pp0_iter2_reg;
            o_1_reg_860_pp0_iter4_reg <= o_1_reg_860_pp0_iter3_reg;
            o_1_reg_860_pp0_iter5_reg <= o_1_reg_860_pp0_iter4_reg;
            o_1_reg_860_pp0_iter6_reg <= o_1_reg_860_pp0_iter5_reg;
            o_1_reg_860_pp0_iter7_reg <= o_1_reg_860_pp0_iter6_reg;
            o_1_reg_860_pp0_iter8_reg <= o_1_reg_860_pp0_iter7_reg;
            o_1_reg_860_pp0_iter9_reg <= o_1_reg_860_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            mul1_i_reg_1050 <= grp_fu_2431_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            mul3_i_reg_1020 <= grp_fu_2443_p_dout0;
            mul6_i_reg_1015 <= grp_fu_2439_p_dout0;
            mul_i_reg_1010  <= grp_fu_2435_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            mul4_i_reg_1025 <= grp_fu_2431_p_dout0;
            mul5_i_reg_1030 <= grp_fu_2435_p_dout0;
            mul7_i_reg_1035 <= grp_fu_2439_p_dout0;
            mul8_i_reg_1040 <= grp_fu_2443_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            mul9_i_reg_1045 <= grp_fu_2431_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            nums_6_reg_887 <= grp_fu_2431_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            nums_6_reg_887_pp0_iter10_reg <= nums_6_reg_887_pp0_iter9_reg;
            nums_6_reg_887_pp0_iter11_reg <= nums_6_reg_887_pp0_iter10_reg;
            nums_6_reg_887_pp0_iter12_reg <= nums_6_reg_887_pp0_iter11_reg;
            nums_6_reg_887_pp0_iter13_reg <= nums_6_reg_887_pp0_iter12_reg;
            nums_6_reg_887_pp0_iter14_reg <= nums_6_reg_887_pp0_iter13_reg;
            nums_6_reg_887_pp0_iter15_reg <= nums_6_reg_887_pp0_iter14_reg;
            nums_6_reg_887_pp0_iter16_reg <= nums_6_reg_887_pp0_iter15_reg;
            nums_6_reg_887_pp0_iter17_reg <= nums_6_reg_887_pp0_iter16_reg;
            nums_6_reg_887_pp0_iter18_reg <= nums_6_reg_887_pp0_iter17_reg;
            nums_6_reg_887_pp0_iter3_reg  <= nums_6_reg_887;
            nums_6_reg_887_pp0_iter4_reg  <= nums_6_reg_887_pp0_iter3_reg;
            nums_6_reg_887_pp0_iter5_reg  <= nums_6_reg_887_pp0_iter4_reg;
            nums_6_reg_887_pp0_iter6_reg  <= nums_6_reg_887_pp0_iter5_reg;
            nums_6_reg_887_pp0_iter7_reg  <= nums_6_reg_887_pp0_iter6_reg;
            nums_6_reg_887_pp0_iter8_reg  <= nums_6_reg_887_pp0_iter7_reg;
            nums_6_reg_887_pp0_iter9_reg  <= nums_6_reg_887_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)))) begin
            reg_609 <= grp_fu_2403_p_dout0;
            reg_615 <= grp_fu_2407_p_dout0;
            reg_621 <= grp_fu_2411_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter26 == 1'b1)))) begin
            reg_627 <= grp_fu_2415_p_dout0;
            reg_634 <= grp_fu_2419_p_dout0;
            reg_641 <= grp_fu_2423_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)))) begin
            reg_648 <= grp_fu_2427_p_dout0;
            reg_655 <= grp_fu_577_p2;
            reg_662 <= grp_fu_581_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            sub204_1_i_reg_1208 <= grp_fu_2407_p_dout0;
            sub204_2_i_reg_1214 <= grp_fu_2411_p_dout0;
            sub7_i_reg_1202 <= grp_fu_2403_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            xL_1_reg_1061 <= grp_fu_2439_p_dout0;
            xL_2_reg_1067 <= grp_fu_2443_p_dout0;
            xL_reg_1055   <= grp_fu_2435_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            yL_1_reg_1080 <= grp_fu_2439_p_dout0;
            yL_2_reg_1087 <= grp_fu_2443_p_dout0;
            yL_reg_1073   <= grp_fu_2435_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            zL_1_reg_1101 <= grp_fu_2435_p_dout0;
            zL_reg_1094   <= grp_fu_2431_p_dout0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln38_reg_867 == 1'd1) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
            ap_condition_exit_pp0_iter0_stage4 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage4 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (icmp_ln38_reg_867_pp0_iter25_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_condition_exit_pp0_iter25_stage1 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter25_stage1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_loop_exit_ready_pp0_iter25_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter26 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to24 = 1'b1;
        end else begin
            ap_idle_pp0_0to24 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter26 == 1'b0))) begin
            ap_idle_pp0_1to26 = 1'b1;
        end else begin
            ap_idle_pp0_1to26 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_o_1 = 4'd0;
        end else begin
            ap_sig_allocacmp_o_1 = o_fu_108;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            env_axesObs_address0 = zext_ln64_9_fu_848_p1;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            env_axesObs_address0 = zext_ln64_8_fu_838_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            env_axesObs_address0 = zext_ln64_5_fu_808_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            env_axesObs_address0 = zext_ln64_3_fu_788_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            env_axesObs_address0 = zext_ln64_1_fu_767_p1;
        end else begin
            env_axesObs_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            env_axesObs_address1 = zext_ln64_7_fu_828_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            env_axesObs_address1 = zext_ln64_6_fu_818_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            env_axesObs_address1 = zext_ln64_4_fu_798_p1;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            env_axesObs_address1 = zext_ln64_2_fu_778_p1;
        end else begin
            env_axesObs_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            env_axesObs_ce0 = 1'b1;
        end else begin
            env_axesObs_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            env_axesObs_ce1 = 1'b1;
        end else begin
            env_axesObs_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            env_axesObs_d0 = H_2_2_reg_958;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            env_axesObs_d0 = H_1_2_reg_933;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            env_axesObs_d0 = H_1_1_reg_927;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            env_axesObs_d0 = H_2_0_reg_946;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            env_axesObs_d0 = H_0_0_reg_896;
        end else begin
            env_axesObs_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            env_axesObs_d1 = H_0_2_reg_908;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            env_axesObs_d1 = H_2_1_reg_952;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            env_axesObs_d1 = H_0_1_reg_902;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            env_axesObs_d1 = H_1_0_reg_921;
        end else begin
            env_axesObs_d1 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            env_axesObs_we0 = 1'b1;
        end else begin
            env_axesObs_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            env_axesObs_we1 = 1'b1;
        end else begin
            env_axesObs_we1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_0_we0 = 1'b1;
        end else begin
            env_pointsObs_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_1_we0 = 1'b1;
        end else begin
            env_pointsObs_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_0_2_we0 = 1'b1;
        end else begin
            env_pointsObs_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_0_we0 = 1'b1;
        end else begin
            env_pointsObs_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_1_we0 = 1'b1;
        end else begin
            env_pointsObs_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_1_2_we0 = 1'b1;
        end else begin
            env_pointsObs_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_0_we0 = 1'b1;
        end else begin
            env_pointsObs_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_1_we0 = 1'b1;
        end else begin
            env_pointsObs_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_2_2_we0 = 1'b1;
        end else begin
            env_pointsObs_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_0_we0 = 1'b1;
        end else begin
            env_pointsObs_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_1_we0 = 1'b1;
        end else begin
            env_pointsObs_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            env_pointsObs_3_2_we0 = 1'b1;
        end else begin
            env_pointsObs_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_4_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_0_we0 = 1'b1;
        end else begin
            env_pointsObs_4_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_4_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_1_we0 = 1'b1;
        end else begin
            env_pointsObs_4_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_4_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            env_pointsObs_4_2_we0 = 1'b1;
        end else begin
            env_pointsObs_4_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_5_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_0_we0 = 1'b1;
        end else begin
            env_pointsObs_5_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_5_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_1_we0 = 1'b1;
        end else begin
            env_pointsObs_5_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_5_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_5_2_we0 = 1'b1;
        end else begin
            env_pointsObs_5_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_6_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_0_we0 = 1'b1;
        end else begin
            env_pointsObs_6_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_6_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_1_we0 = 1'b1;
        end else begin
            env_pointsObs_6_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_6_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_6_2_we0 = 1'b1;
        end else begin
            env_pointsObs_6_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_7_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_0_we0 = 1'b1;
        end else begin
            env_pointsObs_7_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_7_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_1_we0 = 1'b1;
        end else begin
            env_pointsObs_7_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_7_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter25 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            env_pointsObs_7_2_we0 = 1'b1;
        end else begin
            env_pointsObs_7_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_0_ce0 = 1'b1;
        end else begin
            env_pointsObs_8_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_0_we0 = 1'b1;
        end else begin
            env_pointsObs_8_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_1_ce0 = 1'b1;
        end else begin
            env_pointsObs_8_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_1_we0 = 1'b1;
        end else begin
            env_pointsObs_8_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_2_ce0 = 1'b1;
        end else begin
            env_pointsObs_8_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            env_pointsObs_8_2_we0 = 1'b1;
        end else begin
            env_pointsObs_8_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_00001))) begin
            grp_fu_549_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001)))) begin
            grp_fu_549_opcode = 2'd0;
        end else begin
            grp_fu_549_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_549_p0 = add5_i_reg_1184;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_549_p0 = add2_i_reg_1151;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_549_p0 = sub5_i_reg_1133;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_549_p0 = add_i_reg_1115;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_549_p0 = xL_reg_1055;
        end else begin
            grp_fu_549_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_549_p1 = zL_reg_1094_pp0_iter23_reg;
        end else if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_549_p1 = yL_reg_1073_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_549_p1 = H_0_3_reg_914_pp0_iter20_reg;
        end else begin
            grp_fu_549_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_00001))) begin
            grp_fu_553_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001)))) begin
            grp_fu_553_opcode = 2'd0;
        end else begin
            grp_fu_553_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_553_p0 = add158_1_i_reg_1190;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_553_p0 = add67_1_i_reg_1157;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_553_p0 = sub155_1_i_reg_1139;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_553_p0 = add_1_i_reg_1121;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_553_p0 = xL_1_reg_1061;
        end else begin
            grp_fu_553_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_553_p1 = zL_1_reg_1101_pp0_iter23_reg;
        end else if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_553_p1 = yL_1_reg_1080_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_553_p1 = H_1_3_reg_939_pp0_iter20_reg;
        end else begin
            grp_fu_553_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_00001))) begin
            grp_fu_557_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001)))) begin
            grp_fu_557_opcode = 2'd0;
        end else begin
            grp_fu_557_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_557_p0 = add158_2_i_reg_1196;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_557_p0 = add67_2_i_reg_1163;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_557_p0 = sub155_2_i_reg_1145;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_557_p0 = add_2_i_reg_1127;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_557_p0 = xL_2_reg_1067;
        end else begin
            grp_fu_557_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_557_p1 = zL_2_reg_1108_pp0_iter23_reg;
        end else if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_557_p1 = yL_2_reg_1087_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_557_p1 = H_2_3_reg_964_pp0_iter20_reg;
        end else begin
            grp_fu_557_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_561_p0 = sub7_i_reg_1202;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_561_p0 = add5_i_reg_1184;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_561_p0 = add2_i_reg_1151;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_561_p0 = add_i_reg_1115;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_561_p0 = H_0_3_reg_914_pp0_iter20_reg;
        end else begin
            grp_fu_561_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_561_p1 = zL_reg_1094_pp0_iter24_reg;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_561_p1 = zL_reg_1094_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_561_p1 = yL_reg_1073_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_561_p1 = xL_reg_1055;
        end else begin
            grp_fu_561_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_565_p0 = sub204_1_i_reg_1208;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_565_p0 = add158_1_i_reg_1190;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_565_p0 = add67_1_i_reg_1157;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_565_p0 = add_1_i_reg_1121;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_565_p0 = H_1_3_reg_939_pp0_iter20_reg;
        end else begin
            grp_fu_565_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_565_p1 = zL_1_reg_1101_pp0_iter24_reg;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_565_p1 = zL_1_reg_1101_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_565_p1 = yL_1_reg_1080_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_565_p1 = xL_1_reg_1061;
        end else begin
            grp_fu_565_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_569_p0 = sub204_2_i_reg_1214;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_569_p0 = add158_2_i_reg_1196;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_569_p0 = add67_2_i_reg_1163;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_569_p0 = add_2_i_reg_1127;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_569_p0 = H_2_3_reg_964_pp0_iter20_reg;
        end else begin
            grp_fu_569_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_569_p1 = zL_2_reg_1108_pp0_iter24_reg;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_569_p1 = zL_2_reg_1108_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_569_p1 = yL_2_reg_1087_pp0_iter22_reg;
        end else if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_569_p1 = xL_2_reg_1067;
        end else begin
            grp_fu_569_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001))) begin
            grp_fu_573_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)))) begin
            grp_fu_573_opcode = 2'd0;
        end else begin
            grp_fu_573_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_573_p0 = sub7_i_reg_1202;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_573_p0 = sub3_i_reg_1169;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_573_p0 = sub5_i_reg_1133;
        end else begin
            grp_fu_573_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_573_p1 = zL_reg_1094_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_573_p1 = yL_reg_1073_pp0_iter22_reg;
        end else begin
            grp_fu_573_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001))) begin
            grp_fu_577_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)))) begin
            grp_fu_577_opcode = 2'd0;
        end else begin
            grp_fu_577_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_577_p0 = sub204_1_i_reg_1208;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_577_p0 = sub112_1_i_reg_1174;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_577_p0 = sub155_1_i_reg_1139;
        end else begin
            grp_fu_577_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_577_p1 = zL_1_reg_1101_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_577_p1 = yL_1_reg_1080_pp0_iter22_reg;
        end else begin
            grp_fu_577_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001))) begin
            grp_fu_581_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001)))) begin
            grp_fu_581_opcode = 2'd0;
        end else begin
            grp_fu_581_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_581_p0 = sub204_2_i_reg_1214;
        end else if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_581_p0 = sub112_2_i_reg_1179;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_581_p0 = sub155_2_i_reg_1145;
        end else begin
            grp_fu_581_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_581_p1 = zL_2_reg_1108_pp0_iter23_reg;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_581_p1 = yL_2_reg_1087_pp0_iter22_reg;
        end else begin
            grp_fu_581_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_585_p0 = mul8_i_reg_1040;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_585_p0 = H_2_2_reg_958;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_585_p0 = H_1_2_reg_933;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_585_p0 = H_0_1_reg_902;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_585_p0 = conv_i_reg_882;
        end else begin
            grp_fu_585_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_585_p1 = 64'd4602678819172646912;
        end else if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_585_p1 = nums_6_reg_887_pp0_iter18_reg;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_585_p1 = nums_6_reg_887_pp0_iter17_reg;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_585_p1 = 64'd4597094355634707497;
        end else begin
            grp_fu_585_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_590_p0 = mul9_i_reg_1045;
        end else if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_590_p0 = mul4_i_reg_1025;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_590_p0 = mul_i_reg_1010;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_590_p0 = H_1_1_reg_927;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_590_p0 = H_0_0_reg_896;
        end else begin
            grp_fu_590_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_590_p1 = 64'd4602678819172646912;
        end else if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)))) begin
            grp_fu_590_p1 = nums_6_reg_887_pp0_iter17_reg;
        end else begin
            grp_fu_590_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_594_p0 = mul1_i_reg_1050;
        end else if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_594_p0 = mul5_i_reg_1030;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_594_p0 = mul6_i_reg_1015;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_594_p0 = H_2_1_reg_952;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_594_p0 = H_1_0_reg_921;
        end else begin
            grp_fu_594_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1)) | ((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_594_p1 = 64'd4602678819172646912;
        end else if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)))) begin
            grp_fu_594_p1 = nums_6_reg_887_pp0_iter17_reg;
        end else begin
            grp_fu_594_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_598_p0 = mul7_i_reg_1035;
        end else if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_598_p0 = mul3_i_reg_1020;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_598_p0 = H_0_2_reg_908;
        end else if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_598_p0 = H_2_0_reg_946;
        end else begin
            grp_fu_598_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)) | ((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)))) begin
            grp_fu_598_p1 = 64'd4602678819172646912;
        end else if ((((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2)) | ((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3)))) begin
            grp_fu_598_p1 = nums_6_reg_887_pp0_iter17_reg;
        end else begin
            grp_fu_598_p1 = 'bx;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to26 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if (((1'b1 == ap_condition_exit_pp0_iter25_stage1) & (ap_idle_pp0_0to24 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln64_1_fu_772_p2 = (add_ln64_fu_761_p2 + 7'd1);

    assign add_ln64_2_fu_783_p2 = (add_ln64_reg_999 + 7'd2);

    assign add_ln64_3_fu_793_p2 = (add_ln64_reg_999 + 7'd3);

    assign add_ln64_4_fu_803_p2 = (add_ln64_reg_999 + 7'd4);

    assign add_ln64_5_fu_813_p2 = (add_ln64_reg_999 + 7'd5);

    assign add_ln64_6_fu_823_p2 = (add_ln64_reg_999 + 7'd6);

    assign add_ln64_7_fu_833_p2 = (add_ln64_reg_999 + 7'd7);

    assign add_ln64_8_fu_843_p2 = (add_ln64_reg_999 + 7'd8);

    assign add_ln64_fu_761_p2 = (tmp_37_fu_754_p3 + zext_ln64_fu_751_p1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage4;

    assign env_pointsObs_0_0_address0 = zext_ln38_fu_745_p1;

    assign env_pointsObs_0_0_d0 = H_0_3_reg_914;

    assign env_pointsObs_0_1_address0 = zext_ln38_fu_745_p1;

    assign env_pointsObs_0_1_d0 = H_1_3_reg_939;

    assign env_pointsObs_0_2_address0 = zext_ln38_fu_745_p1;

    assign env_pointsObs_0_2_d0 = H_2_3_reg_964;

    assign env_pointsObs_1_0_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_1_0_d0 = reg_609;

    assign env_pointsObs_1_1_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_1_1_d0 = reg_615;

    assign env_pointsObs_1_2_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_1_2_d0 = reg_621;

    assign env_pointsObs_2_0_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_2_0_d0 = reg_627;

    assign env_pointsObs_2_1_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_2_1_d0 = reg_634;

    assign env_pointsObs_2_2_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_2_2_d0 = reg_641;

    assign env_pointsObs_3_0_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_3_0_d0 = reg_648;

    assign env_pointsObs_3_1_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_3_1_d0 = reg_655;

    assign env_pointsObs_3_2_address0 = zext_ln38_reg_971_pp0_iter24_reg;

    assign env_pointsObs_3_2_d0 = reg_662;

    assign env_pointsObs_4_0_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_4_0_d0 = reg_648;

    assign env_pointsObs_4_1_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_4_1_d0 = reg_655;

    assign env_pointsObs_4_2_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_4_2_d0 = reg_662;

    assign env_pointsObs_5_0_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_5_0_d0 = reg_609;

    assign env_pointsObs_5_1_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_5_1_d0 = reg_615;

    assign env_pointsObs_5_2_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_5_2_d0 = reg_621;

    assign env_pointsObs_6_0_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_6_0_d0 = reg_627;

    assign env_pointsObs_6_1_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_6_1_d0 = reg_634;

    assign env_pointsObs_6_2_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_6_2_d0 = reg_641;

    assign env_pointsObs_7_0_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_7_0_d0 = reg_648;

    assign env_pointsObs_7_1_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_7_1_d0 = reg_655;

    assign env_pointsObs_7_2_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_7_2_d0 = reg_662;

    assign env_pointsObs_8_0_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_8_0_d0 = reg_627;

    assign env_pointsObs_8_1_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_8_1_d0 = reg_634;

    assign env_pointsObs_8_2_address0 = zext_ln38_reg_971_pp0_iter25_reg;

    assign env_pointsObs_8_2_d0 = reg_641;

    assign grp_fu_2403_p_ce = 1'b1;

    assign grp_fu_2403_p_din0 = grp_fu_549_p0;

    assign grp_fu_2403_p_din1 = grp_fu_549_p1;

    assign grp_fu_2403_p_opcode = grp_fu_549_opcode;

    assign grp_fu_2407_p_ce = 1'b1;

    assign grp_fu_2407_p_din0 = grp_fu_553_p0;

    assign grp_fu_2407_p_din1 = grp_fu_553_p1;

    assign grp_fu_2407_p_opcode = grp_fu_553_opcode;

    assign grp_fu_2411_p_ce = 1'b1;

    assign grp_fu_2411_p_din0 = grp_fu_557_p0;

    assign grp_fu_2411_p_din1 = grp_fu_557_p1;

    assign grp_fu_2411_p_opcode = grp_fu_557_opcode;

    assign grp_fu_2415_p_ce = 1'b1;

    assign grp_fu_2415_p_din0 = grp_fu_561_p0;

    assign grp_fu_2415_p_din1 = grp_fu_561_p1;

    assign grp_fu_2415_p_opcode = 2'd1;

    assign grp_fu_2419_p_ce = 1'b1;

    assign grp_fu_2419_p_din0 = grp_fu_565_p0;

    assign grp_fu_2419_p_din1 = grp_fu_565_p1;

    assign grp_fu_2419_p_opcode = 2'd1;

    assign grp_fu_2423_p_ce = 1'b1;

    assign grp_fu_2423_p_din0 = grp_fu_569_p0;

    assign grp_fu_2423_p_din1 = grp_fu_569_p1;

    assign grp_fu_2423_p_opcode = 2'd1;

    assign grp_fu_2427_p_ce = 1'b1;

    assign grp_fu_2427_p_din0 = grp_fu_573_p0;

    assign grp_fu_2427_p_din1 = grp_fu_573_p1;

    assign grp_fu_2427_p_opcode = grp_fu_573_opcode;

    assign grp_fu_2431_p_ce = 1'b1;

    assign grp_fu_2431_p_din0 = grp_fu_585_p0;

    assign grp_fu_2431_p_din1 = grp_fu_585_p1;

    assign grp_fu_2435_p_ce = 1'b1;

    assign grp_fu_2435_p_din0 = grp_fu_590_p0;

    assign grp_fu_2435_p_din1 = grp_fu_590_p1;

    assign grp_fu_2439_p_ce = 1'b1;

    assign grp_fu_2439_p_din0 = grp_fu_594_p0;

    assign grp_fu_2439_p_din1 = grp_fu_594_p1;

    assign grp_fu_2443_p_ce = 1'b1;

    assign grp_fu_2443_p_din0 = grp_fu_598_p0;

    assign grp_fu_2443_p_din1 = grp_fu_598_p1;

    assign grp_fu_606_p0 = indvars_iv_next29_i_reg_871;

    assign icmp_ln38_fu_677_p2 = ((ap_sig_allocacmp_o_1 == 4'd8) ? 1'b1 : 1'b0);

    assign indvars_iv_next29_i_fu_683_p2 = (ap_sig_allocacmp_o_1 + 4'd1);

    assign tmp_37_fu_754_p3 = {{o_1_reg_860_pp0_iter18_reg}, {3'd0}};

    assign zext_ln38_fu_745_p1 = o_1_reg_860_pp0_iter18_reg;

    assign zext_ln64_1_fu_767_p1 = add_ln64_fu_761_p2;

    assign zext_ln64_2_fu_778_p1 = add_ln64_1_fu_772_p2;

    assign zext_ln64_3_fu_788_p1 = add_ln64_2_fu_783_p2;

    assign zext_ln64_4_fu_798_p1 = add_ln64_3_fu_793_p2;

    assign zext_ln64_5_fu_808_p1 = add_ln64_4_fu_803_p2;

    assign zext_ln64_6_fu_818_p1 = add_ln64_5_fu_813_p2;

    assign zext_ln64_7_fu_828_p1 = add_ln64_6_fu_823_p2;

    assign zext_ln64_8_fu_838_p1 = add_ln64_7_fu_833_p2;

    assign zext_ln64_9_fu_848_p1 = add_ln64_8_fu_843_p2;

    assign zext_ln64_fu_751_p1 = o_1_reg_860_pp0_iter18_reg;

    always @(posedge ap_clk) begin
        zext_ln38_reg_971[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter19_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter20_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter21_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter22_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter23_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter24_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
        zext_ln38_reg_971_pp0_iter25_reg[63:4] <= 60'b000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_main_Pipeline_VITIS_LOOP_38_1
