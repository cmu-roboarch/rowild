/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_pointsOverlap_double_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    axis_address0,
    axis_ce0,
    axis_q0,
    axis_address1,
    axis_ce1,
    axis_q1,
    axis_offset1,
    ap_return
);

    parameter ap_ST_fsm_pp0_stage0 = 14'd1;
    parameter ap_ST_fsm_pp0_stage1 = 14'd2;
    parameter ap_ST_fsm_pp0_stage2 = 14'd4;
    parameter ap_ST_fsm_pp0_stage3 = 14'd8;
    parameter ap_ST_fsm_pp0_stage4 = 14'd16;
    parameter ap_ST_fsm_pp0_stage5 = 14'd32;
    parameter ap_ST_fsm_pp0_stage6 = 14'd64;
    parameter ap_ST_fsm_pp0_stage7 = 14'd128;
    parameter ap_ST_fsm_pp0_stage8 = 14'd256;
    parameter ap_ST_fsm_pp0_stage9 = 14'd512;
    parameter ap_ST_fsm_pp0_stage10 = 14'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 14'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 14'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 14'd8192;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    output [6:0] axis_address0;
    output axis_ce0;
    input [63:0] axis_q0;
    output [6:0] axis_address1;
    output axis_ce1;
    input [63:0] axis_q1;
    input [1:0] axis_offset1;
    output [0:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[6:0] p1_address0;
    reg p1_ce0;
    reg[6:0] p1_address1;
    reg p1_ce1;
    reg p2_0_0_ce0;
    reg p2_0_1_ce0;
    reg p2_0_2_ce0;
    reg p2_1_0_ce0;
    reg p2_1_1_ce0;
    reg p2_1_2_ce0;
    reg p2_2_0_ce0;
    reg p2_2_1_ce0;
    reg p2_2_2_ce0;
    reg p2_3_0_ce0;
    reg p2_3_1_ce0;
    reg p2_3_2_ce0;
    reg p2_4_0_ce0;
    reg p2_4_1_ce0;
    reg p2_4_2_ce0;
    reg p2_5_0_ce0;
    reg p2_5_1_ce0;
    reg p2_5_2_ce0;
    reg p2_6_0_ce0;
    reg p2_6_1_ce0;
    reg p2_6_2_ce0;
    reg p2_7_0_ce0;
    reg p2_7_1_ce0;
    reg p2_7_2_ce0;
    reg p2_8_0_ce0;
    reg p2_8_1_ce0;
    reg p2_8_2_ce0;
    reg[6:0] axis_address0;
    reg axis_ce0;
    reg axis_ce1;

    (* fsm_encoding = "none" *) reg   [13:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_subdone;
    reg   [63:0] reg_815;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    reg   [63:0] reg_820;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    reg   [63:0] reg_826;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    reg   [63:0] reg_831;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    reg   [63:0] reg_838;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    wire    ap_block_pp0_stage13_11001;
    reg   [63:0] reg_845;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] grp_fu_777_p2;
    reg   [63:0] reg_851;
    wire   [63:0] grp_fu_782_p2;
    reg   [63:0] reg_858;
    reg   [63:0] reg_865;
    reg   [63:0] reg_872;
    reg   [63:0] reg_879;
    reg   [63:0] reg_886;
    reg   [63:0] reg_894;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    reg   [63:0] reg_901;
    reg   [63:0] reg_907;
    reg   [63:0] reg_913;
    wire   [63:0] grp_fu_767_p2;
    reg   [63:0] reg_919;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire   [63:0] p2_offset_cast_fu_930_p1;
    reg   [63:0] p2_offset_cast_reg_3742;
    wire   [6:0] add_ln120_fu_986_p2;
    reg   [6:0] add_ln120_reg_3747;
    wire   [6:0] mul_ln120_fu_996_p2;
    reg   [6:0] mul_ln120_reg_3753;
    wire   [6:0] sub_ln120_2_fu_1012_p2;
    reg   [6:0] sub_ln120_2_reg_3918;
    reg   [63:0] p1_load_reg_3943;
    reg   [63:0] p2_0_0_load_reg_3948;
    reg   [63:0] p2_0_1_load_reg_3953;
    reg   [63:0] p2_0_2_load_reg_3958;
    reg   [63:0] p2_1_0_load_reg_3963;
    reg   [63:0] p2_1_1_load_reg_3968;
    reg   [63:0] p2_1_2_load_reg_3973;
    reg   [63:0] p2_2_0_load_reg_3978;
    reg   [63:0] p2_2_1_load_reg_3983;
    reg   [63:0] p2_2_2_load_reg_3988;
    reg   [63:0] p2_3_0_load_reg_3993;
    reg   [63:0] p2_3_1_load_reg_3998;
    reg   [63:0] p2_3_2_load_reg_4003;
    reg   [63:0] p2_4_0_load_reg_4008;
    reg   [63:0] p2_4_1_load_reg_4013;
    reg   [63:0] p2_4_2_load_reg_4018;
    reg   [63:0] p2_5_0_load_reg_4023;
    reg   [63:0] p2_5_1_load_reg_4028;
    reg   [63:0] p2_5_2_load_reg_4033;
    reg   [63:0] p2_6_0_load_reg_4038;
    reg   [63:0] p2_6_1_load_reg_4043;
    reg   [63:0] p2_6_2_load_reg_4048;
    reg   [63:0] p2_7_0_load_reg_4053;
    reg   [63:0] p2_7_1_load_reg_4058;
    reg   [63:0] p2_7_2_load_reg_4063;
    reg   [63:0] p2_8_0_load_reg_4068;
    reg   [63:0] p2_8_1_load_reg_4073;
    reg   [63:0] axis_load_reg_4093;
    reg   [63:0] axis_load_1_reg_4101;
    reg   [63:0] p1_load_6_reg_4109;
    reg   [63:0] axis_load_2_reg_4124;
    reg   [63:0] p1_load_12_reg_4132;
    reg   [63:0] p1_load_4_reg_4147;
    reg   [63:0] p1_load_7_reg_4162;
    reg   [63:0] p1_load_10_reg_4177;
    reg   [63:0] p1_load_13_reg_4192;
    reg   [63:0] p1_load_2_reg_4207;
    reg   [63:0] p1_load_5_reg_4212;
    wire   [63:0] grp_fu_787_p2;
    reg   [63:0] mul_reg_4227;
    wire   [63:0] grp_fu_791_p2;
    reg   [63:0] mul6_reg_4232;
    wire   [63:0] grp_fu_795_p2;
    reg   [63:0] mul1_reg_4237;
    wire   [63:0] grp_fu_799_p2;
    reg   [63:0] mul2_reg_4242;
    reg   [63:0] p1_load_16_reg_4247;
    reg   [63:0] mul20_1_reg_4262;
    reg   [63:0] mul25_1_reg_4267;
    reg   [63:0] mul20_2_reg_4272;
    reg   [63:0] mul25_2_reg_4277;
    reg   [63:0] p1_load_19_reg_4282;
    reg   [63:0] mul_1_reg_4297;
    reg   [63:0] mul6_1_reg_4302;
    reg   [63:0] mul20_3_reg_4307;
    reg   [63:0] mul25_3_reg_4312;
    reg   [63:0] p1_load_22_reg_4317;
    reg   [63:0] mul20_s_reg_4332;
    reg   [63:0] mul25_s_reg_4337;
    reg   [63:0] mul20_4_reg_4342;
    reg   [63:0] mul25_4_reg_4347;
    reg   [63:0] p1_load_25_reg_4352;
    reg   [63:0] mul20_1_1_reg_4367;
    reg   [63:0] mul25_1_1_reg_4372;
    reg   [63:0] mul20_5_reg_4377;
    reg   [63:0] mul25_5_reg_4382;
    reg   [63:0] p1_load_20_reg_4387;
    reg   [63:0] mul20_2_1_reg_4392;
    reg   [63:0] mul25_2_1_reg_4397;
    reg   [63:0] mul20_6_reg_4402;
    reg   [63:0] mul25_6_reg_4407;
    reg   [63:0] p1_load_26_reg_4412;
    reg   [63:0] mul_2_reg_4422;
    reg   [63:0] mul6_2_reg_4427;
    reg   [63:0] mul20_3_1_reg_4432;
    reg   [63:0] mul25_3_1_reg_4437;
    reg   [63:0] p2_8_2_load_reg_4442;
    reg   [63:0] max1_22_reg_4447;
    wire   [63:0] grp_fu_772_p2;
    reg   [63:0] max2_22_reg_4452;
    reg   [63:0] mul20_8_reg_4457;
    reg   [63:0] mul25_8_reg_4462;
    reg   [63:0] mul20_7_reg_4467;
    reg   [63:0] mul25_7_reg_4472;
    reg   [63:0] n1_3_reg_4477;
    reg   [63:0] n2_3_reg_4482;
    reg   [63:0] mul20_1_2_reg_4487;
    reg   [63:0] mul25_1_2_reg_4492;
    reg   [63:0] n2_6_reg_4497;
    reg   [63:0] mul20_4_1_reg_4502;
    reg   [63:0] mul25_4_1_reg_4507;
    reg   [63:0] mul20_2_2_reg_4512;
    reg   [63:0] mul25_2_2_reg_4517;
    reg   [63:0] n1_9_reg_4522;
    reg   [63:0] n2_9_reg_4527;
    reg   [63:0] mul20_5_1_reg_4532;
    reg   [63:0] mul25_5_1_reg_4537;
    reg   [63:0] mul20_3_2_reg_4542;
    reg   [63:0] mul25_3_2_reg_4547;
    reg   [63:0] n1_26_reg_4552;
    reg   [63:0] n2_26_reg_4557;
    reg   [63:0] mul20_6_1_reg_4562;
    reg   [63:0] mul25_6_1_reg_4567;
    reg   [63:0] mul20_4_2_reg_4572;
    reg   [63:0] mul25_4_2_reg_4577;
    reg   [63:0] n1_29_reg_4582;
    reg   [63:0] n2_29_reg_4587;
    reg   [63:0] mul20_7_1_reg_4592;
    reg   [63:0] mul25_7_1_reg_4597;
    reg   [63:0] mul20_5_2_reg_4602;
    reg   [63:0] mul25_5_2_reg_4607;
    reg   [63:0] n1_32_reg_4612;
    reg   [63:0] n2_32_reg_4617;
    reg   [63:0] mul20_6_2_reg_4622;
    reg   [63:0] mul20_6_2_reg_4622_pp0_iter2_reg;
    reg   [63:0] mul25_6_2_reg_4627;
    reg   [63:0] mul25_6_2_reg_4627_pp0_iter2_reg;
    reg   [63:0] mul20_7_2_reg_4632;
    reg   [63:0] mul20_7_2_reg_4632_pp0_iter2_reg;
    reg   [63:0] mul25_7_2_reg_4637;
    reg   [63:0] mul25_7_2_reg_4637_pp0_iter2_reg;
    reg   [63:0] max1_1_reg_4642;
    reg   [63:0] max2_1_reg_4647;
    reg   [63:0] n1_4_reg_4652;
    reg   [63:0] n2_4_reg_4657;
    reg   [63:0] n1_7_reg_4662;
    reg   [63:0] n2_7_reg_4667;
    reg   [63:0] n1_24_reg_4672;
    reg   [63:0] n2_24_reg_4677;
    reg   [63:0] n1_35_reg_4682;
    reg   [63:0] n2_35_reg_4687;
    reg   [63:0] n1_27_reg_4692;
    reg   [63:0] n2_27_reg_4697;
    reg   [63:0] n1_30_reg_4702;
    reg   [63:0] n2_30_reg_4707;
    reg   [63:0] n1_33_reg_4712;
    reg   [63:0] n2_33_reg_4717;
    wire   [63:0] max1_fu_1387_p3;
    reg   [63:0] max1_reg_4722;
    wire   [63:0] min1_11_fu_1401_p3;
    reg   [63:0] min1_11_reg_4729;
    wire   [0:0] and_ln135_fu_1481_p2;
    reg   [0:0] and_ln135_reg_4736;
    wire   [0:0] grp_fu_811_p2;
    reg   [0:0] tmp_93_reg_4742;
    wire   [63:0] max2_fu_1491_p3;
    reg   [63:0] max2_reg_4747;
    wire   [63:0] min2_11_fu_1505_p3;
    reg   [63:0] min2_11_reg_4754;
    reg   [63:0] n2_25_reg_4761;
    reg   [63:0] n1_36_reg_4770;
    wire   [63:0] max1_15_fu_1596_p3;
    reg   [63:0] max1_15_reg_4775;
    wire   [63:0] min1_12_fu_1650_p3;
    reg   [63:0] min1_12_reg_4782;
    wire   [0:0] or_ln135_17_fu_1704_p2;
    reg   [0:0] or_ln135_17_reg_4789;
    wire   [63:0] max2_15_fu_1740_p3;
    reg   [63:0] max2_15_reg_4794;
    wire   [63:0] min2_12_fu_1793_p3;
    reg   [63:0] min2_12_reg_4801;
    wire   [63:0] max1_16_fu_1883_p3;
    reg   [63:0] max1_16_reg_4808;
    wire   [63:0] min1_13_fu_1937_p3;
    reg   [63:0] min1_13_reg_4815;
    wire   [0:0] or_ln135_19_fu_1991_p2;
    reg   [0:0] or_ln135_19_reg_4822;
    wire   [63:0] max2_16_fu_2027_p3;
    reg   [63:0] max2_16_reg_4827;
    wire   [63:0] min2_13_fu_2080_p3;
    reg   [63:0] min2_13_reg_4834;
    wire   [63:0] max1_17_fu_2170_p3;
    reg   [63:0] max1_17_reg_4841;
    wire   [63:0] min1_14_fu_2224_p3;
    reg   [63:0] min1_14_reg_4848;
    wire   [0:0] or_ln135_21_fu_2277_p2;
    reg   [0:0] or_ln135_21_reg_4855;
    wire   [63:0] max2_17_fu_2313_p3;
    reg   [63:0] max2_17_reg_4860;
    wire   [63:0] min2_14_fu_2365_p3;
    reg   [63:0] min2_14_reg_4867;
    wire   [63:0] max1_18_fu_2454_p3;
    reg   [63:0] max1_18_reg_4874;
    wire   [63:0] min1_15_fu_2508_p3;
    reg   [63:0] min1_15_reg_4881;
    wire   [0:0] or_ln135_23_fu_2562_p2;
    reg   [0:0] or_ln135_23_reg_4888;
    wire   [63:0] max2_18_fu_2598_p3;
    reg   [63:0] max2_18_reg_4893;
    reg   [63:0] n2_37_reg_4900;
    wire   [63:0] min2_15_fu_2651_p3;
    reg   [63:0] min2_15_reg_4909;
    wire   [63:0] max1_19_fu_2741_p3;
    reg   [63:0] max1_19_reg_4916;
    wire   [63:0] min1_16_fu_2795_p3;
    reg   [63:0] min1_16_reg_4923;
    wire   [0:0] or_ln135_25_fu_2849_p2;
    reg   [0:0] or_ln135_25_reg_4930;
    wire   [63:0] max2_19_fu_2885_p3;
    reg   [63:0] max2_19_reg_4935;
    wire   [63:0] min2_16_fu_2938_p3;
    reg   [63:0] min2_16_reg_4942;
    wire   [63:0] max1_20_fu_3028_p3;
    reg   [63:0] max1_20_reg_4949;
    wire   [63:0] min1_17_fu_3082_p3;
    reg   [63:0] min1_17_reg_4956;
    wire   [0:0] or_ln135_27_fu_3136_p2;
    reg   [0:0] or_ln135_27_reg_4963;
    wire   [63:0] max2_20_fu_3172_p3;
    reg   [63:0] max2_20_reg_4968;
    wire   [63:0] min2_17_fu_3225_p3;
    reg   [63:0] min2_17_reg_4975;
    wire   [63:0] max1_21_fu_3315_p3;
    reg   [63:0] max1_21_reg_4982;
    wire   [63:0] min1_18_fu_3369_p3;
    reg   [63:0] min1_18_reg_4989;
    wire   [63:0] max2_21_fu_3458_p3;
    reg   [63:0] max2_21_reg_4997;
    wire   [63:0] min2_18_fu_3511_p3;
    reg   [63:0] min2_18_reg_5005;
    wire   [0:0] grp_fu_807_p2;
    reg   [0:0] tmp_169_reg_5012;
    reg   [0:0] tmp_171_reg_5017;
    reg   [0:0] tmp_172_reg_5022;
    reg   [0:0] tmp_173_reg_5027;
    wire   [0:0] and_ln139_5_fu_3587_p2;
    reg   [0:0] and_ln139_5_reg_5032;
    wire   [0:0] and_ln139_8_fu_3634_p2;
    reg   [0:0] and_ln139_8_reg_5037;
    wire   [0:0] and_ln140_7_fu_3685_p2;
    reg   [0:0] and_ln140_7_reg_5043;
    wire   [0:0] and_ln140_fu_3707_p2;
    reg   [0:0] and_ln140_reg_5048;
    reg   [0:0] tmp_167_reg_5053;
    wire   [0:0] or_ln140_5_fu_3723_p2;
    reg   [0:0] or_ln140_5_reg_5058;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage3_subdone;
    wire   [63:0] zext_ln120_14_fu_1002_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln120_10_fu_1017_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln120_11_fu_1028_p1;
    wire   [63:0] zext_ln129_fu_1038_p1;
    wire   [63:0] zext_ln129_26_fu_1048_p1;
    wire   [63:0] zext_ln120_12_fu_1058_p1;
    wire    ap_block_pp0_stage2;
    wire   [63:0] zext_ln129_29_fu_1068_p1;
    wire   [63:0] zext_ln129_32_fu_1078_p1;
    wire   [63:0] zext_ln120_15_fu_1088_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln129_24_fu_1098_p1;
    wire   [63:0] zext_ln129_27_fu_1108_p1;
    wire    ap_block_pp0_stage4;
    wire   [63:0] zext_ln129_35_fu_1118_p1;
    wire   [63:0] zext_ln129_30_fu_1128_p1;
    wire    ap_block_pp0_stage5;
    wire   [63:0] zext_ln129_38_fu_1138_p1;
    wire   [63:0] zext_ln129_33_fu_1148_p1;
    wire    ap_block_pp0_stage6;
    wire   [63:0] zext_ln129_41_fu_1158_p1;
    wire   [63:0] zext_ln120_16_fu_1168_p1;
    wire    ap_block_pp0_stage7;
    wire   [63:0] zext_ln129_25_fu_1178_p1;
    wire   [63:0] zext_ln129_36_fu_1188_p1;
    wire    ap_block_pp0_stage8;
    wire   [63:0] zext_ln129_44_fu_1198_p1;
    wire   [63:0] zext_ln129_28_fu_1208_p1;
    wire    ap_block_pp0_stage9;
    wire   [63:0] zext_ln129_39_fu_1218_p1;
    wire   [63:0] zext_ln129_31_fu_1228_p1;
    wire    ap_block_pp0_stage10;
    wire   [63:0] zext_ln129_42_fu_1238_p1;
    wire   [63:0] zext_ln129_34_fu_1248_p1;
    wire    ap_block_pp0_stage11;
    wire   [63:0] zext_ln129_45_fu_1258_p1;
    wire   [63:0] zext_ln129_37_fu_1268_p1;
    wire    ap_block_pp0_stage12;
    wire   [63:0] zext_ln129_40_fu_1278_p1;
    wire   [63:0] zext_ln129_43_fu_1288_p1;
    wire    ap_block_pp0_stage13;
    wire   [63:0] zext_ln129_46_fu_1298_p1;
    reg   [63:0] grp_fu_767_p0;
    reg   [63:0] grp_fu_767_p1;
    reg   [63:0] grp_fu_772_p0;
    reg   [63:0] grp_fu_772_p1;
    reg   [63:0] grp_fu_777_p0;
    reg   [63:0] grp_fu_777_p1;
    reg   [63:0] grp_fu_782_p0;
    reg   [63:0] grp_fu_782_p1;
    reg   [63:0] grp_fu_787_p0;
    reg   [63:0] grp_fu_787_p1;
    reg   [63:0] grp_fu_791_p0;
    reg   [63:0] grp_fu_791_p1;
    reg   [63:0] grp_fu_795_p0;
    reg   [63:0] grp_fu_795_p1;
    reg   [63:0] grp_fu_799_p0;
    reg   [63:0] grp_fu_799_p1;
    reg   [63:0] grp_fu_803_p0;
    reg   [63:0] grp_fu_803_p1;
    reg   [63:0] grp_fu_807_p0;
    reg   [63:0] grp_fu_807_p1;
    reg   [63:0] grp_fu_811_p0;
    reg   [63:0] grp_fu_811_p1;
    wire   [4:0] tmp_fu_964_p3;
    wire   [5:0] zext_ln120_9_fu_972_p1;
    wire   [5:0] zext_ln120_fu_960_p1;
    wire   [5:0] sub_ln120_fu_976_p2;
    wire  signed [6:0] sext_ln120_fu_982_p1;
    wire   [6:0] axis_offset1_cast3_fu_926_p1;
    wire   [1:0] mul_ln120_fu_996_p0;
    wire   [5:0] mul_ln120_fu_996_p1;
    wire   [6:0] shl_ln120_fu_1007_p2;
    wire   [6:0] add_ln120_5_fu_1022_p2;
    wire   [6:0] add_ln129_fu_1033_p2;
    wire   [6:0] add_ln129_26_fu_1043_p2;
    wire   [6:0] add_ln120_6_fu_1053_p2;
    wire   [6:0] add_ln129_29_fu_1063_p2;
    wire   [6:0] add_ln129_32_fu_1073_p2;
    wire   [6:0] add_ln120_7_fu_1083_p2;
    wire   [6:0] add_ln129_24_fu_1093_p2;
    wire   [6:0] add_ln129_27_fu_1103_p2;
    wire   [6:0] add_ln129_35_fu_1113_p2;
    wire   [6:0] add_ln129_30_fu_1123_p2;
    wire   [6:0] add_ln129_38_fu_1133_p2;
    wire   [6:0] add_ln129_33_fu_1143_p2;
    wire   [6:0] add_ln129_41_fu_1153_p2;
    wire   [6:0] add_ln120_8_fu_1163_p2;
    wire   [6:0] add_ln129_25_fu_1173_p2;
    wire   [6:0] add_ln129_36_fu_1183_p2;
    wire   [6:0] add_ln129_44_fu_1193_p2;
    wire   [6:0] add_ln129_28_fu_1203_p2;
    wire   [6:0] add_ln129_39_fu_1213_p2;
    wire   [6:0] add_ln129_31_fu_1223_p2;
    wire   [6:0] add_ln129_42_fu_1233_p2;
    wire   [6:0] add_ln129_34_fu_1243_p2;
    wire   [6:0] add_ln129_45_fu_1253_p2;
    wire   [6:0] add_ln129_37_fu_1263_p2;
    wire   [6:0] add_ln129_40_fu_1273_p2;
    wire   [6:0] add_ln129_43_fu_1283_p2;
    wire   [6:0] add_ln129_46_fu_1293_p2;
    wire   [63:0] bitcast_ln133_fu_1303_p1;
    wire   [63:0] bitcast_ln133_16_fu_1321_p1;
    wire   [10:0] tmp_s_fu_1307_p4;
    wire   [51:0] trunc_ln133_fu_1317_p1;
    wire   [0:0] icmp_ln133_32_fu_1345_p2;
    wire   [0:0] icmp_ln133_fu_1339_p2;
    wire   [10:0] tmp_88_fu_1325_p4;
    wire   [51:0] trunc_ln133_16_fu_1335_p1;
    wire   [0:0] icmp_ln133_34_fu_1363_p2;
    wire   [0:0] icmp_ln133_33_fu_1357_p2;
    wire   [0:0] or_ln133_fu_1351_p2;
    wire   [0:0] or_ln133_16_fu_1369_p2;
    wire   [0:0] and_ln133_fu_1375_p2;
    wire   [0:0] grp_fu_803_p2;
    wire   [0:0] and_ln133_16_fu_1381_p2;
    wire   [0:0] and_ln134_fu_1395_p2;
    wire   [63:0] bitcast_ln135_fu_1409_p1;
    wire   [63:0] bitcast_ln135_16_fu_1427_p1;
    wire   [10:0] tmp_91_fu_1413_p4;
    wire   [51:0] trunc_ln135_fu_1423_p1;
    wire   [0:0] icmp_ln135_32_fu_1451_p2;
    wire   [0:0] icmp_ln135_fu_1445_p2;
    wire   [10:0] tmp_92_fu_1431_p4;
    wire   [51:0] trunc_ln135_16_fu_1441_p1;
    wire   [0:0] icmp_ln135_34_fu_1469_p2;
    wire   [0:0] icmp_ln135_33_fu_1463_p2;
    wire   [0:0] or_ln135_fu_1457_p2;
    wire   [0:0] or_ln135_16_fu_1475_p2;
    wire   [0:0] and_ln135_16_fu_1487_p2;
    wire   [0:0] and_ln136_fu_1500_p2;
    wire   [63:0] bitcast_ln133_17_fu_1513_p1;
    wire   [63:0] bitcast_ln133_18_fu_1531_p1;
    wire   [10:0] tmp_95_fu_1517_p4;
    wire   [51:0] trunc_ln133_17_fu_1527_p1;
    wire   [0:0] icmp_ln133_36_fu_1554_p2;
    wire   [0:0] icmp_ln133_35_fu_1548_p2;
    wire   [10:0] tmp_96_fu_1534_p4;
    wire   [51:0] trunc_ln133_18_fu_1544_p1;
    wire   [0:0] icmp_ln133_38_fu_1572_p2;
    wire   [0:0] icmp_ln133_37_fu_1566_p2;
    wire   [0:0] or_ln133_17_fu_1560_p2;
    wire   [0:0] or_ln133_18_fu_1578_p2;
    wire   [0:0] and_ln133_17_fu_1584_p2;
    wire   [0:0] and_ln133_18_fu_1590_p2;
    wire   [63:0] bitcast_ln134_fu_1603_p1;
    wire   [10:0] tmp_98_fu_1606_p4;
    wire   [51:0] trunc_ln134_fu_1616_p1;
    wire   [0:0] icmp_ln134_14_fu_1626_p2;
    wire   [0:0] icmp_ln134_fu_1620_p2;
    wire   [0:0] or_ln134_fu_1632_p2;
    wire   [0:0] and_ln134_15_fu_1638_p2;
    wire   [0:0] and_ln134_16_fu_1644_p2;
    wire   [63:0] bitcast_ln135_17_fu_1657_p1;
    wire   [63:0] bitcast_ln135_18_fu_1675_p1;
    wire   [10:0] tmp_100_fu_1661_p4;
    wire   [51:0] trunc_ln135_17_fu_1671_p1;
    wire   [0:0] icmp_ln135_36_fu_1698_p2;
    wire   [0:0] icmp_ln135_35_fu_1692_p2;
    wire   [10:0] tmp_101_fu_1678_p4;
    wire   [51:0] trunc_ln135_18_fu_1688_p1;
    wire   [0:0] icmp_ln135_38_fu_1716_p2;
    wire   [0:0] icmp_ln135_37_fu_1710_p2;
    wire   [0:0] or_ln135_18_fu_1722_p2;
    wire   [0:0] and_ln135_17_fu_1728_p2;
    wire   [0:0] and_ln135_18_fu_1734_p2;
    wire   [63:0] bitcast_ln136_fu_1747_p1;
    wire   [10:0] tmp_103_fu_1750_p4;
    wire   [51:0] trunc_ln136_fu_1760_p1;
    wire   [0:0] icmp_ln136_14_fu_1770_p2;
    wire   [0:0] icmp_ln136_fu_1764_p2;
    wire   [0:0] or_ln136_fu_1776_p2;
    wire   [0:0] and_ln136_15_fu_1782_p2;
    wire   [0:0] and_ln136_16_fu_1787_p2;
    wire   [63:0] bitcast_ln133_19_fu_1800_p1;
    wire   [63:0] bitcast_ln133_20_fu_1818_p1;
    wire   [10:0] tmp_105_fu_1804_p4;
    wire   [51:0] trunc_ln133_19_fu_1814_p1;
    wire   [0:0] icmp_ln133_40_fu_1841_p2;
    wire   [0:0] icmp_ln133_39_fu_1835_p2;
    wire   [10:0] tmp_106_fu_1821_p4;
    wire   [51:0] trunc_ln133_20_fu_1831_p1;
    wire   [0:0] icmp_ln133_42_fu_1859_p2;
    wire   [0:0] icmp_ln133_41_fu_1853_p2;
    wire   [0:0] or_ln133_19_fu_1847_p2;
    wire   [0:0] or_ln133_20_fu_1865_p2;
    wire   [0:0] and_ln133_19_fu_1871_p2;
    wire   [0:0] and_ln133_20_fu_1877_p2;
    wire   [63:0] bitcast_ln134_7_fu_1890_p1;
    wire   [10:0] tmp_108_fu_1893_p4;
    wire   [51:0] trunc_ln134_7_fu_1903_p1;
    wire   [0:0] icmp_ln134_16_fu_1913_p2;
    wire   [0:0] icmp_ln134_15_fu_1907_p2;
    wire   [0:0] or_ln134_7_fu_1919_p2;
    wire   [0:0] and_ln134_17_fu_1925_p2;
    wire   [0:0] and_ln134_18_fu_1931_p2;
    wire   [63:0] bitcast_ln135_19_fu_1944_p1;
    wire   [63:0] bitcast_ln135_20_fu_1962_p1;
    wire   [10:0] tmp_110_fu_1948_p4;
    wire   [51:0] trunc_ln135_19_fu_1958_p1;
    wire   [0:0] icmp_ln135_40_fu_1985_p2;
    wire   [0:0] icmp_ln135_39_fu_1979_p2;
    wire   [10:0] tmp_111_fu_1965_p4;
    wire   [51:0] trunc_ln135_20_fu_1975_p1;
    wire   [0:0] icmp_ln135_42_fu_2003_p2;
    wire   [0:0] icmp_ln135_41_fu_1997_p2;
    wire   [0:0] or_ln135_20_fu_2009_p2;
    wire   [0:0] and_ln135_19_fu_2015_p2;
    wire   [0:0] and_ln135_20_fu_2021_p2;
    wire   [63:0] bitcast_ln136_7_fu_2034_p1;
    wire   [10:0] tmp_113_fu_2037_p4;
    wire   [51:0] trunc_ln136_7_fu_2047_p1;
    wire   [0:0] icmp_ln136_16_fu_2057_p2;
    wire   [0:0] icmp_ln136_15_fu_2051_p2;
    wire   [0:0] or_ln136_7_fu_2063_p2;
    wire   [0:0] and_ln136_17_fu_2069_p2;
    wire   [0:0] and_ln136_18_fu_2074_p2;
    wire   [63:0] bitcast_ln133_21_fu_2087_p1;
    wire   [63:0] bitcast_ln133_22_fu_2105_p1;
    wire   [10:0] tmp_115_fu_2091_p4;
    wire   [51:0] trunc_ln133_21_fu_2101_p1;
    wire   [0:0] icmp_ln133_44_fu_2128_p2;
    wire   [0:0] icmp_ln133_43_fu_2122_p2;
    wire   [10:0] tmp_116_fu_2108_p4;
    wire   [51:0] trunc_ln133_22_fu_2118_p1;
    wire   [0:0] icmp_ln133_46_fu_2146_p2;
    wire   [0:0] icmp_ln133_45_fu_2140_p2;
    wire   [0:0] or_ln133_21_fu_2134_p2;
    wire   [0:0] or_ln133_22_fu_2152_p2;
    wire   [0:0] and_ln133_21_fu_2158_p2;
    wire   [0:0] and_ln133_22_fu_2164_p2;
    wire   [63:0] bitcast_ln134_8_fu_2177_p1;
    wire   [10:0] tmp_118_fu_2180_p4;
    wire   [51:0] trunc_ln134_8_fu_2190_p1;
    wire   [0:0] icmp_ln134_18_fu_2200_p2;
    wire   [0:0] icmp_ln134_17_fu_2194_p2;
    wire   [0:0] or_ln134_8_fu_2206_p2;
    wire   [0:0] and_ln134_19_fu_2212_p2;
    wire   [0:0] and_ln134_20_fu_2218_p2;
    wire   [63:0] bitcast_ln135_21_fu_2231_p1;
    wire   [63:0] bitcast_ln135_22_fu_2248_p1;
    wire   [10:0] tmp_120_fu_2234_p4;
    wire   [51:0] trunc_ln135_21_fu_2244_p1;
    wire   [0:0] icmp_ln135_44_fu_2271_p2;
    wire   [0:0] icmp_ln135_43_fu_2265_p2;
    wire   [10:0] tmp_121_fu_2251_p4;
    wire   [51:0] trunc_ln135_22_fu_2261_p1;
    wire   [0:0] icmp_ln135_46_fu_2289_p2;
    wire   [0:0] icmp_ln135_45_fu_2283_p2;
    wire   [0:0] or_ln135_22_fu_2295_p2;
    wire   [0:0] and_ln135_21_fu_2301_p2;
    wire   [0:0] and_ln135_22_fu_2307_p2;
    wire   [63:0] bitcast_ln136_8_fu_2319_p1;
    wire   [10:0] tmp_123_fu_2322_p4;
    wire   [51:0] trunc_ln136_8_fu_2332_p1;
    wire   [0:0] icmp_ln136_18_fu_2342_p2;
    wire   [0:0] icmp_ln136_17_fu_2336_p2;
    wire   [0:0] or_ln136_8_fu_2348_p2;
    wire   [0:0] and_ln136_19_fu_2354_p2;
    wire   [0:0] and_ln136_20_fu_2359_p2;
    wire   [63:0] bitcast_ln133_23_fu_2371_p1;
    wire   [63:0] bitcast_ln133_24_fu_2389_p1;
    wire   [10:0] tmp_125_fu_2375_p4;
    wire   [51:0] trunc_ln133_23_fu_2385_p1;
    wire   [0:0] icmp_ln133_48_fu_2412_p2;
    wire   [0:0] icmp_ln133_47_fu_2406_p2;
    wire   [10:0] tmp_126_fu_2392_p4;
    wire   [51:0] trunc_ln133_24_fu_2402_p1;
    wire   [0:0] icmp_ln133_50_fu_2430_p2;
    wire   [0:0] icmp_ln133_49_fu_2424_p2;
    wire   [0:0] or_ln133_23_fu_2418_p2;
    wire   [0:0] or_ln133_24_fu_2436_p2;
    wire   [0:0] and_ln133_23_fu_2442_p2;
    wire   [0:0] and_ln133_24_fu_2448_p2;
    wire   [63:0] bitcast_ln134_9_fu_2461_p1;
    wire   [10:0] tmp_128_fu_2464_p4;
    wire   [51:0] trunc_ln134_9_fu_2474_p1;
    wire   [0:0] icmp_ln134_20_fu_2484_p2;
    wire   [0:0] icmp_ln134_19_fu_2478_p2;
    wire   [0:0] or_ln134_9_fu_2490_p2;
    wire   [0:0] and_ln134_21_fu_2496_p2;
    wire   [0:0] and_ln134_22_fu_2502_p2;
    wire   [63:0] bitcast_ln135_23_fu_2515_p1;
    wire   [63:0] bitcast_ln135_24_fu_2533_p1;
    wire   [10:0] tmp_130_fu_2519_p4;
    wire   [51:0] trunc_ln135_23_fu_2529_p1;
    wire   [0:0] icmp_ln135_48_fu_2556_p2;
    wire   [0:0] icmp_ln135_47_fu_2550_p2;
    wire   [10:0] tmp_131_fu_2536_p4;
    wire   [51:0] trunc_ln135_24_fu_2546_p1;
    wire   [0:0] icmp_ln135_50_fu_2574_p2;
    wire   [0:0] icmp_ln135_49_fu_2568_p2;
    wire   [0:0] or_ln135_24_fu_2580_p2;
    wire   [0:0] and_ln135_23_fu_2586_p2;
    wire   [0:0] and_ln135_24_fu_2592_p2;
    wire   [63:0] bitcast_ln136_9_fu_2605_p1;
    wire   [10:0] tmp_133_fu_2608_p4;
    wire   [51:0] trunc_ln136_9_fu_2618_p1;
    wire   [0:0] icmp_ln136_20_fu_2628_p2;
    wire   [0:0] icmp_ln136_19_fu_2622_p2;
    wire   [0:0] or_ln136_9_fu_2634_p2;
    wire   [0:0] and_ln136_21_fu_2640_p2;
    wire   [0:0] and_ln136_22_fu_2645_p2;
    wire   [63:0] bitcast_ln133_25_fu_2658_p1;
    wire   [63:0] bitcast_ln133_26_fu_2676_p1;
    wire   [10:0] tmp_135_fu_2662_p4;
    wire   [51:0] trunc_ln133_25_fu_2672_p1;
    wire   [0:0] icmp_ln133_52_fu_2699_p2;
    wire   [0:0] icmp_ln133_51_fu_2693_p2;
    wire   [10:0] tmp_136_fu_2679_p4;
    wire   [51:0] trunc_ln133_26_fu_2689_p1;
    wire   [0:0] icmp_ln133_54_fu_2717_p2;
    wire   [0:0] icmp_ln133_53_fu_2711_p2;
    wire   [0:0] or_ln133_25_fu_2705_p2;
    wire   [0:0] or_ln133_26_fu_2723_p2;
    wire   [0:0] and_ln133_25_fu_2729_p2;
    wire   [0:0] and_ln133_26_fu_2735_p2;
    wire   [63:0] bitcast_ln134_10_fu_2748_p1;
    wire   [10:0] tmp_138_fu_2751_p4;
    wire   [51:0] trunc_ln134_10_fu_2761_p1;
    wire   [0:0] icmp_ln134_22_fu_2771_p2;
    wire   [0:0] icmp_ln134_21_fu_2765_p2;
    wire   [0:0] or_ln134_10_fu_2777_p2;
    wire   [0:0] and_ln134_23_fu_2783_p2;
    wire   [0:0] and_ln134_24_fu_2789_p2;
    wire   [63:0] bitcast_ln135_25_fu_2802_p1;
    wire   [63:0] bitcast_ln135_26_fu_2820_p1;
    wire   [10:0] tmp_140_fu_2806_p4;
    wire   [51:0] trunc_ln135_25_fu_2816_p1;
    wire   [0:0] icmp_ln135_52_fu_2843_p2;
    wire   [0:0] icmp_ln135_51_fu_2837_p2;
    wire   [10:0] tmp_141_fu_2823_p4;
    wire   [51:0] trunc_ln135_26_fu_2833_p1;
    wire   [0:0] icmp_ln135_54_fu_2861_p2;
    wire   [0:0] icmp_ln135_53_fu_2855_p2;
    wire   [0:0] or_ln135_26_fu_2867_p2;
    wire   [0:0] and_ln135_25_fu_2873_p2;
    wire   [0:0] and_ln135_26_fu_2879_p2;
    wire   [63:0] bitcast_ln136_10_fu_2892_p1;
    wire   [10:0] tmp_143_fu_2895_p4;
    wire   [51:0] trunc_ln136_10_fu_2905_p1;
    wire   [0:0] icmp_ln136_22_fu_2915_p2;
    wire   [0:0] icmp_ln136_21_fu_2909_p2;
    wire   [0:0] or_ln136_10_fu_2921_p2;
    wire   [0:0] and_ln136_23_fu_2927_p2;
    wire   [0:0] and_ln136_24_fu_2932_p2;
    wire   [63:0] bitcast_ln133_27_fu_2945_p1;
    wire   [63:0] bitcast_ln133_28_fu_2963_p1;
    wire   [10:0] tmp_145_fu_2949_p4;
    wire   [51:0] trunc_ln133_27_fu_2959_p1;
    wire   [0:0] icmp_ln133_56_fu_2986_p2;
    wire   [0:0] icmp_ln133_55_fu_2980_p2;
    wire   [10:0] tmp_146_fu_2966_p4;
    wire   [51:0] trunc_ln133_28_fu_2976_p1;
    wire   [0:0] icmp_ln133_58_fu_3004_p2;
    wire   [0:0] icmp_ln133_57_fu_2998_p2;
    wire   [0:0] or_ln133_27_fu_2992_p2;
    wire   [0:0] or_ln133_28_fu_3010_p2;
    wire   [0:0] and_ln133_27_fu_3016_p2;
    wire   [0:0] and_ln133_28_fu_3022_p2;
    wire   [63:0] bitcast_ln134_11_fu_3035_p1;
    wire   [10:0] tmp_148_fu_3038_p4;
    wire   [51:0] trunc_ln134_11_fu_3048_p1;
    wire   [0:0] icmp_ln134_24_fu_3058_p2;
    wire   [0:0] icmp_ln134_23_fu_3052_p2;
    wire   [0:0] or_ln134_11_fu_3064_p2;
    wire   [0:0] and_ln134_25_fu_3070_p2;
    wire   [0:0] and_ln134_26_fu_3076_p2;
    wire   [63:0] bitcast_ln135_27_fu_3089_p1;
    wire   [63:0] bitcast_ln135_28_fu_3107_p1;
    wire   [10:0] tmp_150_fu_3093_p4;
    wire   [51:0] trunc_ln135_27_fu_3103_p1;
    wire   [0:0] icmp_ln135_56_fu_3130_p2;
    wire   [0:0] icmp_ln135_55_fu_3124_p2;
    wire   [10:0] tmp_151_fu_3110_p4;
    wire   [51:0] trunc_ln135_28_fu_3120_p1;
    wire   [0:0] icmp_ln135_58_fu_3148_p2;
    wire   [0:0] icmp_ln135_57_fu_3142_p2;
    wire   [0:0] or_ln135_28_fu_3154_p2;
    wire   [0:0] and_ln135_27_fu_3160_p2;
    wire   [0:0] and_ln135_28_fu_3166_p2;
    wire   [63:0] bitcast_ln136_11_fu_3179_p1;
    wire   [10:0] tmp_153_fu_3182_p4;
    wire   [51:0] trunc_ln136_11_fu_3192_p1;
    wire   [0:0] icmp_ln136_24_fu_3202_p2;
    wire   [0:0] icmp_ln136_23_fu_3196_p2;
    wire   [0:0] or_ln136_11_fu_3208_p2;
    wire   [0:0] and_ln136_25_fu_3214_p2;
    wire   [0:0] and_ln136_26_fu_3219_p2;
    wire   [63:0] bitcast_ln133_29_fu_3232_p1;
    wire   [63:0] bitcast_ln133_30_fu_3250_p1;
    wire   [10:0] tmp_155_fu_3236_p4;
    wire   [51:0] trunc_ln133_29_fu_3246_p1;
    wire   [0:0] icmp_ln133_60_fu_3273_p2;
    wire   [0:0] icmp_ln133_59_fu_3267_p2;
    wire   [10:0] tmp_156_fu_3253_p4;
    wire   [51:0] trunc_ln133_30_fu_3263_p1;
    wire   [0:0] icmp_ln133_62_fu_3291_p2;
    wire   [0:0] icmp_ln133_61_fu_3285_p2;
    wire   [0:0] or_ln133_29_fu_3279_p2;
    wire   [0:0] or_ln133_30_fu_3297_p2;
    wire   [0:0] and_ln133_29_fu_3303_p2;
    wire   [0:0] and_ln133_30_fu_3309_p2;
    wire   [63:0] bitcast_ln134_12_fu_3322_p1;
    wire   [10:0] tmp_158_fu_3325_p4;
    wire   [51:0] trunc_ln134_12_fu_3335_p1;
    wire   [0:0] icmp_ln134_26_fu_3345_p2;
    wire   [0:0] icmp_ln134_25_fu_3339_p2;
    wire   [0:0] or_ln134_12_fu_3351_p2;
    wire   [0:0] and_ln134_27_fu_3357_p2;
    wire   [0:0] and_ln134_28_fu_3363_p2;
    wire   [63:0] bitcast_ln135_29_fu_3376_p1;
    wire   [63:0] bitcast_ln135_30_fu_3393_p1;
    wire   [10:0] tmp_160_fu_3379_p4;
    wire   [51:0] trunc_ln135_29_fu_3389_p1;
    wire   [0:0] icmp_ln135_60_fu_3416_p2;
    wire   [0:0] icmp_ln135_59_fu_3410_p2;
    wire   [10:0] tmp_161_fu_3396_p4;
    wire   [51:0] trunc_ln135_30_fu_3406_p1;
    wire   [0:0] icmp_ln135_62_fu_3434_p2;
    wire   [0:0] icmp_ln135_61_fu_3428_p2;
    wire   [0:0] or_ln135_29_fu_3422_p2;
    wire   [0:0] or_ln135_30_fu_3440_p2;
    wire   [0:0] and_ln135_29_fu_3446_p2;
    wire   [0:0] and_ln135_30_fu_3452_p2;
    wire   [63:0] bitcast_ln136_12_fu_3464_p1;
    wire   [10:0] tmp_163_fu_3467_p4;
    wire   [51:0] trunc_ln136_12_fu_3477_p1;
    wire   [0:0] icmp_ln136_26_fu_3487_p2;
    wire   [0:0] icmp_ln136_25_fu_3481_p2;
    wire   [0:0] or_ln136_12_fu_3493_p2;
    wire   [0:0] and_ln136_27_fu_3499_p2;
    wire   [0:0] and_ln136_28_fu_3505_p2;
    wire   [63:0] bitcast_ln139_fu_3517_p1;
    wire   [63:0] bitcast_ln139_3_fu_3534_p1;
    wire   [10:0] tmp_165_fu_3520_p4;
    wire   [51:0] trunc_ln139_fu_3530_p1;
    wire   [0:0] icmp_ln139_6_fu_3557_p2;
    wire   [0:0] icmp_ln139_fu_3551_p2;
    wire   [10:0] tmp_166_fu_3537_p4;
    wire   [51:0] trunc_ln139_3_fu_3547_p1;
    wire   [0:0] icmp_ln139_8_fu_3575_p2;
    wire   [0:0] icmp_ln139_7_fu_3569_p2;
    wire   [0:0] or_ln139_fu_3563_p2;
    wire   [0:0] or_ln139_3_fu_3581_p2;
    wire   [63:0] bitcast_ln139_4_fu_3593_p1;
    wire   [10:0] tmp_168_fu_3596_p4;
    wire   [51:0] trunc_ln139_4_fu_3606_p1;
    wire   [0:0] icmp_ln139_10_fu_3616_p2;
    wire   [0:0] icmp_ln139_9_fu_3610_p2;
    wire   [0:0] or_ln139_4_fu_3622_p2;
    wire   [0:0] and_ln139_7_fu_3628_p2;
    wire   [63:0] bitcast_ln140_fu_3639_p1;
    wire   [10:0] tmp_170_fu_3642_p4;
    wire   [51:0] trunc_ln140_fu_3652_p1;
    wire   [0:0] icmp_ln140_2_fu_3662_p2;
    wire   [0:0] icmp_ln140_fu_3656_p2;
    wire   [0:0] or_ln140_4_fu_3668_p2;
    wire   [0:0] and_ln140_5_fu_3674_p2;
    wire   [0:0] and_ln140_8_fu_3691_p2;
    wire   [0:0] and_ln141_fu_3696_p2;
    wire   [0:0] and_ln140_6_fu_3680_p2;
    wire   [0:0] or_ln140_fu_3701_p2;
    wire   [0:0] and_ln142_2_fu_3713_p2;
    wire   [0:0] and_ln142_fu_3718_p2;
    wire   [0:0] and_ln139_6_fu_3728_p2;
    wire   [0:0] and_ln139_fu_3732_p2;
    reg   [4:0] grp_fu_803_opcode;
    wire    ap_block_pp0_stage6_00001;
    wire    ap_block_pp0_stage7_00001;
    wire    ap_block_pp0_stage8_00001;
    wire    ap_block_pp0_stage9_00001;
    wire    ap_block_pp0_stage10_00001;
    wire    ap_block_pp0_stage11_00001;
    wire    ap_block_pp0_stage12_00001;
    wire    ap_block_pp0_stage13_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage5_00001;
    reg   [4:0] grp_fu_807_opcode;
    reg   [4:0] grp_fu_811_opcode;
    reg   [13:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to4;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    reg    ap_idle_pp0_0to3;
    reg    ap_reset_idle_pp0;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_enable_pp0;
    wire   [6:0] mul_ln120_fu_996_p00;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 14'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
    end

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1171 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_767_p0),
        .din1(grp_fu_767_p1),
        .ce(1'b1),
        .dout(grp_fu_767_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1172 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_772_p0),
        .din1(grp_fu_772_p1),
        .ce(1'b1),
        .dout(grp_fu_772_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1173 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_777_p0),
        .din1(grp_fu_777_p1),
        .ce(1'b1),
        .dout(grp_fu_777_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1174 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_782_p0),
        .din1(grp_fu_782_p1),
        .ce(1'b1),
        .dout(grp_fu_782_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1175 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_787_p0),
        .din1(grp_fu_787_p1),
        .ce(1'b1),
        .dout(grp_fu_787_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1176 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_791_p0),
        .din1(grp_fu_791_p1),
        .ce(1'b1),
        .dout(grp_fu_791_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1177 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_795_p0),
        .din1(grp_fu_795_p1),
        .ce(1'b1),
        .dout(grp_fu_795_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U1178 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_799_p0),
        .din1(grp_fu_799_p1),
        .ce(1'b1),
        .dout(grp_fu_799_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1179 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_803_p0),
        .din1(grp_fu_803_p1),
        .ce(1'b1),
        .opcode(grp_fu_803_opcode),
        .dout(grp_fu_803_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1180 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_807_p0),
        .din1(grp_fu_807_p1),
        .ce(1'b1),
        .opcode(grp_fu_807_opcode),
        .dout(grp_fu_807_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_x_U1181 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_811_p0),
        .din1(grp_fu_811_p1),
        .ce(1'b1),
        .opcode(grp_fu_811_opcode),
        .dout(grp_fu_811_p2)
    );

    main_mul_2ns_6ns_7_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(2),
        .din1_WIDTH(6),
        .dout_WIDTH(7)
    ) mul_2ns_6ns_7_1_1_U1182 (
        .din0(mul_ln120_fu_996_p0),
        .din1(mul_ln120_fu_996_p1),
        .dout(mul_ln120_fu_996_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                ap_enable_reg_pp0_iter4 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                reg_831 <= p1_q0;
            end else if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                reg_831 <= p1_q1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13_11001) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                reg_838 <= p1_q0;
            end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                reg_838 <= p1_q1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            reg_845 <= p1_q0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            reg_845 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            add_ln120_reg_3747 <= add_ln120_fu_986_p2;
            min2_14_reg_4867 <= min2_14_fu_2365_p3;
            mul_ln120_reg_3753 <= mul_ln120_fu_996_p2;
            p2_offset_cast_reg_3742[2 : 0] <= p2_offset_cast_fu_930_p1[2 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            and_ln135_reg_4736 <= and_ln135_fu_1481_p2;
            max1_reg_4722 <= max1_fu_1387_p3;
            min1_11_reg_4729 <= min1_11_fu_1401_p3;
            mul20_6_2_reg_4622_pp0_iter2_reg <= mul20_6_2_reg_4622;
            mul25_6_2_reg_4627_pp0_iter2_reg <= mul25_6_2_reg_4627;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            and_ln139_5_reg_5032 <= and_ln139_5_fu_3587_p2;
            and_ln139_8_reg_5037 <= and_ln139_8_fu_3634_p2;
            and_ln140_7_reg_5043 <= and_ln140_7_fu_3685_p2;
            and_ln140_reg_5048 <= and_ln140_fu_3707_p2;
            max1_18_reg_4874 <= max1_18_fu_2454_p3;
            max2_18_reg_4893 <= max2_18_fu_2598_p3;
            min1_15_reg_4881 <= min1_15_fu_2508_p3;
            or_ln135_23_reg_4888 <= or_ln135_23_fu_2562_p2;
            p2_0_0_load_reg_3948 <= p2_0_0_q0;
            p2_0_1_load_reg_3953 <= p2_0_1_q0;
            p2_0_2_load_reg_3958 <= p2_0_2_q0;
            p2_1_0_load_reg_3963 <= p2_1_0_q0;
            p2_1_1_load_reg_3968 <= p2_1_1_q0;
            p2_1_2_load_reg_3973 <= p2_1_2_q0;
            p2_2_0_load_reg_3978 <= p2_2_0_q0;
            p2_2_1_load_reg_3983 <= p2_2_1_q0;
            p2_2_2_load_reg_3988 <= p2_2_2_q0;
            p2_3_0_load_reg_3993 <= p2_3_0_q0;
            p2_3_1_load_reg_3998 <= p2_3_1_q0;
            p2_3_2_load_reg_4003 <= p2_3_2_q0;
            p2_4_0_load_reg_4008 <= p2_4_0_q0;
            p2_4_1_load_reg_4013 <= p2_4_1_q0;
            p2_4_2_load_reg_4018 <= p2_4_2_q0;
            p2_5_0_load_reg_4023 <= p2_5_0_q0;
            p2_5_1_load_reg_4028 <= p2_5_1_q0;
            p2_5_2_load_reg_4033 <= p2_5_2_q0;
            p2_6_0_load_reg_4038 <= p2_6_0_q0;
            p2_6_1_load_reg_4043 <= p2_6_1_q0;
            p2_6_2_load_reg_4048 <= p2_6_2_q0;
            p2_7_0_load_reg_4053 <= p2_7_0_q0;
            p2_7_1_load_reg_4058 <= p2_7_1_q0;
            p2_7_2_load_reg_4063 <= p2_7_2_q0;
            p2_8_0_load_reg_4068 <= p2_8_0_q0;
            p2_8_1_load_reg_4073 <= p2_8_1_q0;
            p2_8_2_load_reg_4442 <= p2_8_2_q0;
            sub_ln120_2_reg_3918 <= sub_ln120_2_fu_1012_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            axis_load_1_reg_4101 <= axis_q0;
            axis_load_reg_4093   <= axis_q1;
            p1_load_6_reg_4109   <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            axis_load_2_reg_4124 <= axis_q0;
            p1_load_12_reg_4132  <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            max1_15_reg_4775 <= max1_15_fu_1596_p3;
            max2_15_reg_4794 <= max2_15_fu_1740_p3;
            min1_12_reg_4782 <= min1_12_fu_1650_p3;
            or_ln135_17_reg_4789 <= or_ln135_17_fu_1704_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            max1_16_reg_4808 <= max1_16_fu_1883_p3;
            max2_16_reg_4827 <= max2_16_fu_2027_p3;
            min1_13_reg_4815 <= min1_13_fu_1937_p3;
            or_ln135_19_reg_4822 <= or_ln135_19_fu_1991_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            max1_17_reg_4841 <= max1_17_fu_2170_p3;
            max2_17_reg_4860 <= max2_17_fu_2313_p3;
            min1_14_reg_4848 <= min1_14_fu_2224_p3;
            or_ln135_21_reg_4855 <= or_ln135_21_fu_2277_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            max1_19_reg_4916 <= max1_19_fu_2741_p3;
            max2_19_reg_4935 <= max2_19_fu_2885_p3;
            min1_16_reg_4923 <= min1_16_fu_2795_p3;
            or_ln135_25_reg_4930 <= or_ln135_25_fu_2849_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            max1_1_reg_4642 <= grp_fu_767_p2;
            max2_1_reg_4647 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            max1_20_reg_4949 <= max1_20_fu_3028_p3;
            max2_20_reg_4968 <= max2_20_fu_3172_p3;
            min1_17_reg_4956 <= min1_17_fu_3082_p3;
            or_ln135_27_reg_4963 <= or_ln135_27_fu_3136_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            max1_21_reg_4982 <= max1_21_fu_3315_p3;
            max2_reg_4747 <= max2_fu_1491_p3;
            min1_18_reg_4989 <= min1_18_fu_3369_p3;
            min2_11_reg_4754 <= min2_11_fu_1505_p3;
            mul20_7_2_reg_4632_pp0_iter2_reg <= mul20_7_2_reg_4632;
            mul25_7_2_reg_4637_pp0_iter2_reg <= mul25_7_2_reg_4637;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            max1_22_reg_4447 <= grp_fu_767_p2;
            max2_22_reg_4452 <= grp_fu_772_p2;
            mul20_7_reg_4467 <= grp_fu_795_p2;
            mul20_8_reg_4457 <= grp_fu_787_p2;
            mul25_7_reg_4472 <= grp_fu_799_p2;
            mul25_8_reg_4462 <= grp_fu_791_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            max2_21_reg_4997 <= max2_21_fu_3458_p3;
            min2_12_reg_4801 <= min2_12_fu_1793_p3;
            min2_18_reg_5005 <= min2_18_fu_3511_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            min2_13_reg_4834 <= min2_13_fu_2080_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            min2_15_reg_4909 <= min2_15_fu_2651_p3;
            or_ln140_5_reg_5058 <= or_ln140_5_fu_3723_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            min2_16_reg_4942 <= min2_16_fu_2938_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            min2_17_reg_4975 <= min2_17_fu_3225_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            mul1_reg_4237 <= grp_fu_795_p2;
            mul2_reg_4242 <= grp_fu_799_p2;
            mul6_reg_4232 <= grp_fu_791_p2;
            mul_reg_4227 <= grp_fu_787_p2;
            p1_load_16_reg_4247 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            mul20_1_1_reg_4367 <= grp_fu_787_p2;
            mul20_5_reg_4377 <= grp_fu_795_p2;
            mul25_1_1_reg_4372 <= grp_fu_791_p2;
            mul25_5_reg_4382 <= grp_fu_799_p2;
            p1_load_20_reg_4387 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            mul20_1_2_reg_4487 <= grp_fu_787_p2;
            mul20_4_1_reg_4502 <= grp_fu_795_p2;
            mul25_1_2_reg_4492 <= grp_fu_791_p2;
            mul25_4_1_reg_4507 <= grp_fu_799_p2;
            n1_3_reg_4477 <= grp_fu_767_p2;
            n2_3_reg_4482 <= grp_fu_772_p2;
            n2_6_reg_4497 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            mul20_1_reg_4262 <= grp_fu_787_p2;
            mul20_2_reg_4272 <= grp_fu_795_p2;
            mul25_1_reg_4267 <= grp_fu_791_p2;
            mul25_2_reg_4277 <= grp_fu_799_p2;
            p1_load_19_reg_4282 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            mul20_2_1_reg_4392 <= grp_fu_787_p2;
            mul20_6_reg_4402 <= grp_fu_795_p2;
            mul25_2_1_reg_4397 <= grp_fu_791_p2;
            mul25_6_reg_4407 <= grp_fu_799_p2;
            p1_load_26_reg_4412 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul20_2_2_reg_4512 <= grp_fu_787_p2;
            mul20_5_1_reg_4532 <= grp_fu_795_p2;
            mul25_2_2_reg_4517 <= grp_fu_791_p2;
            mul25_5_1_reg_4537 <= grp_fu_799_p2;
            n1_9_reg_4522 <= grp_fu_767_p2;
            n2_9_reg_4527 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            mul20_3_1_reg_4432 <= grp_fu_795_p2;
            mul25_3_1_reg_4437 <= grp_fu_799_p2;
            mul6_2_reg_4427 <= grp_fu_791_p2;
            mul_2_reg_4422 <= grp_fu_787_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            mul20_3_2_reg_4542 <= grp_fu_787_p2;
            mul20_6_1_reg_4562 <= grp_fu_795_p2;
            mul25_3_2_reg_4547 <= grp_fu_791_p2;
            mul25_6_1_reg_4567 <= grp_fu_799_p2;
            n1_26_reg_4552 <= grp_fu_767_p2;
            n2_26_reg_4557 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            mul20_3_reg_4307 <= grp_fu_795_p2;
            mul25_3_reg_4312 <= grp_fu_799_p2;
            mul6_1_reg_4302 <= grp_fu_791_p2;
            mul_1_reg_4297 <= grp_fu_787_p2;
            p1_load_22_reg_4317 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            mul20_4_2_reg_4572 <= grp_fu_787_p2;
            mul20_7_1_reg_4592 <= grp_fu_795_p2;
            mul25_4_2_reg_4577 <= grp_fu_791_p2;
            mul25_7_1_reg_4597 <= grp_fu_799_p2;
            n1_29_reg_4582 <= grp_fu_767_p2;
            n2_29_reg_4587 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            mul20_4_reg_4342 <= grp_fu_795_p2;
            mul20_s_reg_4332 <= grp_fu_787_p2;
            mul25_4_reg_4347 <= grp_fu_799_p2;
            mul25_s_reg_4337 <= grp_fu_791_p2;
            p1_load_25_reg_4352 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            mul20_5_2_reg_4602 <= grp_fu_787_p2;
            mul20_6_2_reg_4622 <= grp_fu_795_p2;
            mul25_5_2_reg_4607 <= grp_fu_791_p2;
            mul25_6_2_reg_4627 <= grp_fu_799_p2;
            n1_32_reg_4612 <= grp_fu_767_p2;
            n2_32_reg_4617 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            mul20_7_2_reg_4632 <= grp_fu_787_p2;
            mul25_7_2_reg_4637 <= grp_fu_791_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            n1_24_reg_4672 <= grp_fu_767_p2;
            n1_35_reg_4682 <= grp_fu_777_p2;
            n2_24_reg_4677 <= grp_fu_772_p2;
            n2_35_reg_4687 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            n1_27_reg_4692 <= grp_fu_767_p2;
            n2_27_reg_4697 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            n1_30_reg_4702 <= grp_fu_767_p2;
            n2_30_reg_4707 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            n1_33_reg_4712 <= grp_fu_767_p2;
            n2_33_reg_4717 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            n1_36_reg_4770 <= grp_fu_777_p2;
            n2_25_reg_4761 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            n1_4_reg_4652 <= grp_fu_767_p2;
            n1_7_reg_4662 <= grp_fu_777_p2;
            n2_4_reg_4657 <= grp_fu_772_p2;
            n2_7_reg_4667 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            n2_37_reg_4900 <= grp_fu_772_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            p1_load_10_reg_4177 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            p1_load_13_reg_4192 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            p1_load_2_reg_4207 <= p1_q0;
            p1_load_5_reg_4212 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            p1_load_4_reg_4147 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            p1_load_7_reg_4162 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            p1_load_reg_3943 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            reg_815 <= p1_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_820 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_826 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            reg_851 <= grp_fu_777_p2;
            reg_858 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            reg_865 <= grp_fu_777_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)))) begin
            reg_872 <= grp_fu_777_p2;
            reg_879 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_886 <= grp_fu_777_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            reg_894 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_901 <= grp_fu_777_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_907 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_913 <= grp_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_919 <= grp_fu_767_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            tmp_167_reg_5053 <= grp_fu_807_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            tmp_169_reg_5012 <= grp_fu_807_p2;
            tmp_171_reg_5017 <= grp_fu_811_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            tmp_172_reg_5022 <= grp_fu_807_p2;
            tmp_173_reg_5027 <= grp_fu_811_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            tmp_93_reg_4742 <= grp_fu_811_p2;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to3 = 1'b1;
        end else begin
            ap_idle_pp0_0to3 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to4 = 1'b1;
        end else begin
            ap_idle_pp0_1to4 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0_0to3 == 1'b1) & (ap_start == 1'b0))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                axis_address0 = zext_ln120_12_fu_1058_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                axis_address0 = zext_ln120_11_fu_1028_p1;
            end else begin
                axis_address0 = 'bx;
            end
        end else begin
            axis_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            axis_ce0 = 1'b1;
        end else begin
            axis_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            axis_ce1 = 1'b1;
        end else begin
            axis_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_767_p0 = n1_36_reg_4770;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_767_p0 = n1_24_reg_4672;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_767_p0 = n1_32_reg_4612;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_767_p0 = n1_29_reg_4582;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_767_p0 = n1_26_reg_4552;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_767_p0 = n1_9_reg_4522;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_767_p0 = n1_3_reg_4477;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_767_p0 = max1_22_reg_4447;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_767_p0 = mul20_6_reg_4402;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_767_p0 = mul20_5_reg_4377;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_767_p0 = mul20_4_reg_4342;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_767_p0 = mul20_3_reg_4307;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_767_p0 = mul20_1_reg_4262;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_767_p0 = mul_reg_4227;
        end else begin
            grp_fu_767_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_767_p1 = mul20_7_2_reg_4632_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_767_p1 = mul20_3_2_reg_4542;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_767_p1 = mul20_6_1_reg_4562;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_767_p1 = mul20_5_1_reg_4532;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_767_p1 = mul20_4_1_reg_4502;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_767_p1 = mul20_3_1_reg_4432;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_767_p1 = mul20_1_1_reg_4367;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_767_p1 = mul_1_reg_4297;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_767_p1 = 64'd0;
        end else begin
            grp_fu_767_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_772_p0 = reg_894;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_772_p0 = n2_24_reg_4677;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_772_p0 = n2_32_reg_4617;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_772_p0 = n2_29_reg_4587;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_772_p0 = n2_26_reg_4557;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_772_p0 = n2_9_reg_4527;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_772_p0 = n2_3_reg_4482;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_772_p0 = max2_22_reg_4452;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_772_p0 = mul25_6_reg_4407;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_772_p0 = mul25_5_reg_4382;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_772_p0 = mul25_4_reg_4347;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_772_p0 = mul25_3_reg_4312;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_772_p0 = mul25_1_reg_4267;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_772_p0 = mul6_reg_4232;
        end else begin
            grp_fu_772_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_772_p1 = mul25_7_2_reg_4637_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_772_p1 = mul25_3_2_reg_4547;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_772_p1 = mul25_6_1_reg_4567;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_772_p1 = mul25_5_1_reg_4537;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_772_p1 = mul25_4_1_reg_4507;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_772_p1 = mul25_3_1_reg_4437;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_772_p1 = mul25_1_1_reg_4372;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_772_p1 = mul6_1_reg_4302;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_772_p1 = 64'd0;
        end else begin
            grp_fu_772_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_777_p0 = n1_33_reg_4712;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_777_p0 = n1_30_reg_4702;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_777_p0 = n1_27_reg_4692;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_777_p0 = n1_35_reg_4682;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_777_p0 = n1_7_reg_4662;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_777_p0 = n1_4_reg_4652;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_777_p0 = reg_872;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_777_p0 = max1_1_reg_4642;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_777_p0 = mul20_7_reg_4467;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_777_p0 = reg_865;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_777_p0 = reg_851;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_777_p0 = mul20_2_reg_4272;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_777_p0 = mul1_reg_4237;
        end else begin
            grp_fu_777_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_777_p1 = mul20_6_2_reg_4622_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_777_p1 = mul20_5_2_reg_4602;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_777_p1 = mul20_4_2_reg_4572;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_777_p1 = mul20_7_1_reg_4592;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_777_p1 = mul20_2_2_reg_4512;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_777_p1 = mul20_1_2_reg_4487;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_777_p1 = mul20_8_reg_4457;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_777_p1 = mul_2_reg_4422;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_777_p1 = mul20_2_1_reg_4392;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_777_p1 = mul20_s_reg_4332;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_777_p1 = 64'd0;
        end else begin
            grp_fu_777_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_782_p0 = n2_33_reg_4717;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_782_p0 = n2_30_reg_4707;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_782_p0 = n2_27_reg_4697;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_782_p0 = n2_35_reg_4687;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_782_p0 = n2_7_reg_4667;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_782_p0 = n2_4_reg_4657;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_782_p0 = reg_879;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_782_p0 = max2_1_reg_4647;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_782_p0 = mul25_7_reg_4472;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_782_p0 = n2_6_reg_4497;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_782_p0 = reg_858;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_782_p0 = mul25_2_reg_4277;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_782_p0 = mul2_reg_4242;
        end else begin
            grp_fu_782_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_782_p1 = mul25_6_2_reg_4627_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_782_p1 = mul25_5_2_reg_4607;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_782_p1 = mul25_4_2_reg_4577;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_782_p1 = mul25_7_1_reg_4597;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_782_p1 = mul25_2_2_reg_4517;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_782_p1 = mul25_1_2_reg_4492;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_782_p1 = mul25_8_reg_4462;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_782_p1 = mul6_2_reg_4427;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_782_p1 = mul25_2_1_reg_4397;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_782_p1 = mul25_s_reg_4337;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_782_p1 = 64'd0;
        end else begin
            grp_fu_782_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_787_p0 = p1_load_26_reg_4412;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_787_p0 = p1_load_20_reg_4387;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_787_p0 = reg_838;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_787_p0 = reg_831;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_787_p0 = reg_820;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_787_p0 = p1_load_5_reg_4212;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_787_p0 = p1_load_2_reg_4207;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_787_p0 = p1_load_10_reg_4177;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_787_p0 = p1_load_7_reg_4162;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_787_p0 = p1_load_4_reg_4147;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_787_p0 = reg_826;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_787_p0 = p1_load_6_reg_4109;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_787_p0 = p1_load_reg_3943;
        end else begin
            grp_fu_787_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_787_p1 = axis_load_2_reg_4124;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_787_p1 = axis_load_1_reg_4101;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_787_p1 = axis_load_reg_4093;
        end else begin
            grp_fu_787_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_791_p0 = p2_8_2_load_reg_4442;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_791_p0 = p2_6_2_load_reg_4048;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_791_p0 = p2_5_2_load_reg_4033;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_791_p0 = p2_4_2_load_reg_4018;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_791_p0 = p2_3_2_load_reg_4003;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_791_p0 = p2_2_2_load_reg_3988;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_791_p0 = p2_1_2_load_reg_3973;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_791_p0 = p2_0_2_load_reg_3958;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_791_p0 = p2_3_1_load_reg_3998;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_791_p0 = p2_2_1_load_reg_3983;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_791_p0 = p2_1_1_load_reg_3968;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_791_p0 = p2_0_1_load_reg_3953;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_791_p0 = p2_2_0_load_reg_3978;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_791_p0 = p2_0_0_load_reg_3948;
        end else begin
            grp_fu_791_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_791_p1 = axis_load_2_reg_4124;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_791_p1 = axis_load_1_reg_4101;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_791_p1 = axis_load_reg_4093;
        end else begin
            grp_fu_791_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_795_p0 = p1_load_25_reg_4352;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_795_p0 = p1_load_22_reg_4317;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_795_p0 = p1_load_19_reg_4282;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_795_p0 = p1_load_16_reg_4247;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_795_p0 = p1_load_13_reg_4192;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_795_p0 = reg_845;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_795_p0 = reg_838;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_795_p0 = reg_831;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_795_p0 = p1_load_12_reg_4132;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_795_p0 = reg_820;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_795_p0 = reg_815;
        end else begin
            grp_fu_795_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_795_p1 = axis_load_2_reg_4124;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_795_p1 = axis_load_1_reg_4101;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_795_p1 = axis_load_reg_4093;
        end else begin
            grp_fu_795_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_799_p0 = p2_7_2_load_reg_4063;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_799_p0 = p2_8_1_load_reg_4073;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_799_p0 = p2_7_1_load_reg_4058;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_799_p0 = p2_6_1_load_reg_4043;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_799_p0 = p2_5_1_load_reg_4028;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_799_p0 = p2_8_0_load_reg_4068;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_799_p0 = p2_4_1_load_reg_4013;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_799_p0 = p2_7_0_load_reg_4053;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_799_p0 = p2_6_0_load_reg_4038;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_799_p0 = p2_5_0_load_reg_4023;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_799_p0 = p2_4_0_load_reg_4008;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_799_p0 = p2_3_0_load_reg_3993;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_799_p0 = p2_1_0_load_reg_3963;
        end else begin
            grp_fu_799_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_799_p1 = axis_load_2_reg_4124;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_799_p1 = axis_load_1_reg_4101;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_799_p1 = axis_load_reg_4093;
        end else begin
            grp_fu_799_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_803_opcode = 5'd4;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_803_opcode = 5'd2;
        end else begin
            grp_fu_803_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_803_p0 = reg_865;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_803_p0 = reg_858;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_803_p0 = reg_851;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_803_p0 = n2_25_reg_4761;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_803_p0 = reg_919;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_803_p0 = reg_913;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_803_p0 = reg_886;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_803_p0 = reg_907;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_803_p0 = reg_901;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_803_p0 = reg_879;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_803_p0 = reg_872;
        end else begin
            grp_fu_803_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_803_p1 = min2_16_reg_4942;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_803_p1 = max1_19_reg_4916;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_803_p1 = min2_15_reg_4909;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_803_p1 = max1_18_reg_4874;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_803_p1 = min2_14_reg_4867;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_803_p1 = max1_17_reg_4841;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_803_p1 = min2_13_reg_4834;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_803_p1 = max1_16_reg_4808;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_803_p1 = min2_12_reg_4801;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_803_p1 = max1_15_reg_4775;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_803_p1 = min2_11_reg_4754;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_803_p1 = max1_reg_4722;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_803_p1 = reg_894;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_803_p1 = reg_886;
        end else begin
            grp_fu_803_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_807_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_807_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_807_opcode = 5'd2;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_807_opcode = 5'd4;
        end else begin
            grp_fu_807_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_807_p0 = min1_18_reg_4989;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_807_p0 = max1_21_reg_4982;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_807_p0 = n2_37_reg_4900;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_807_p0 = reg_865;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_807_p0 = reg_851;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_807_p0 = reg_919;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_807_p0 = reg_886;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_807_p0 = reg_901;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_807_p0 = reg_872;
        end else begin
            grp_fu_807_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_807_p1 = max2_21_reg_4997;
        end else if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_807_p1 = min2_18_reg_5005;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_807_p1 = max2_20_reg_4968;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_807_p1 = max1_20_reg_4949;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_807_p1 = min1_16_reg_4923;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_807_p1 = min1_15_reg_4881;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_807_p1 = min1_14_reg_4848;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_807_p1 = min1_13_reg_4815;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_807_p1 = min1_12_reg_4782;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_807_p1 = min1_11_reg_4729;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_807_p1 = reg_886;
        end else begin
            grp_fu_807_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_811_opcode = 5'd3;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_811_opcode = 5'd5;
        end else if ((((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_811_opcode = 5'd4;
        end else if ((((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_811_opcode = 5'd2;
        end else begin
            grp_fu_811_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_811_p0 = min2_18_reg_5005;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_811_p0 = max2_21_reg_4997;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_811_p0 = min1_18_reg_4989;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_811_p0 = n2_37_reg_4900;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_811_p0 = reg_919;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_811_p0 = reg_858;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_811_p0 = n2_25_reg_4761;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_811_p0 = reg_913;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_811_p0 = reg_907;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_811_p0 = reg_879;
        end else begin
            grp_fu_811_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_811_p1 = min1_18_reg_4989;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            grp_fu_811_p1 = max1_21_reg_4982;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            grp_fu_811_p1 = max2_21_reg_4997;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_811_p1 = min2_17_reg_4975;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            grp_fu_811_p1 = min1_17_reg_4956;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_811_p1 = max2_19_reg_4935;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_811_p1 = max2_18_reg_4893;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_811_p1 = max2_17_reg_4860;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            grp_fu_811_p1 = max2_16_reg_4827;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            grp_fu_811_p1 = max2_15_reg_4794;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_811_p1 = max2_fu_1491_p3;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_811_p1 = reg_894;
        end else begin
            grp_fu_811_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address0 = zext_ln129_43_fu_1288_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address0 = zext_ln129_37_fu_1268_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address0 = zext_ln129_34_fu_1248_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address0 = zext_ln129_31_fu_1228_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address0 = zext_ln129_28_fu_1208_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address0 = zext_ln129_36_fu_1188_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address0 = zext_ln120_16_fu_1168_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address0 = zext_ln129_33_fu_1148_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address0 = zext_ln129_30_fu_1128_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address0 = zext_ln129_27_fu_1108_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address0 = zext_ln120_15_fu_1088_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address0 = zext_ln129_29_fu_1068_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address0 = zext_ln129_26_fu_1048_p1;
            end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                p1_address0 = zext_ln120_14_fu_1002_p1;
            end else begin
                p1_address0 = 'bx;
            end
        end else begin
            p1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage13) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                p1_address1 = zext_ln129_46_fu_1298_p1;
            end else if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                p1_address1 = zext_ln129_40_fu_1278_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                p1_address1 = zext_ln129_45_fu_1258_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                p1_address1 = zext_ln129_42_fu_1238_p1;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                p1_address1 = zext_ln129_39_fu_1218_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                p1_address1 = zext_ln129_44_fu_1198_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                p1_address1 = zext_ln129_25_fu_1178_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                p1_address1 = zext_ln129_41_fu_1158_p1;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                p1_address1 = zext_ln129_38_fu_1138_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                p1_address1 = zext_ln129_35_fu_1118_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                p1_address1 = zext_ln129_24_fu_1098_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                p1_address1 = zext_ln129_32_fu_1078_p1;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                p1_address1 = zext_ln129_fu_1038_p1;
            end else begin
                p1_address1 = 'bx;
            end
        end else begin
            p1_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            p1_ce0 = 1'b1;
        end else begin
            p1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage10_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            p1_ce1 = 1'b1;
        end else begin
            p1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_0_ce0 = 1'b1;
        end else begin
            p2_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_1_ce0 = 1'b1;
        end else begin
            p2_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_0_2_ce0 = 1'b1;
        end else begin
            p2_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_0_ce0 = 1'b1;
        end else begin
            p2_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_1_ce0 = 1'b1;
        end else begin
            p2_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_1_2_ce0 = 1'b1;
        end else begin
            p2_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_0_ce0 = 1'b1;
        end else begin
            p2_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_1_ce0 = 1'b1;
        end else begin
            p2_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_2_2_ce0 = 1'b1;
        end else begin
            p2_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_0_ce0 = 1'b1;
        end else begin
            p2_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_1_ce0 = 1'b1;
        end else begin
            p2_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_3_2_ce0 = 1'b1;
        end else begin
            p2_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_0_ce0 = 1'b1;
        end else begin
            p2_4_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_1_ce0 = 1'b1;
        end else begin
            p2_4_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_4_2_ce0 = 1'b1;
        end else begin
            p2_4_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_0_ce0 = 1'b1;
        end else begin
            p2_5_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_1_ce0 = 1'b1;
        end else begin
            p2_5_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_5_2_ce0 = 1'b1;
        end else begin
            p2_5_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_0_ce0 = 1'b1;
        end else begin
            p2_6_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_1_ce0 = 1'b1;
        end else begin
            p2_6_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_6_2_ce0 = 1'b1;
        end else begin
            p2_6_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_0_ce0 = 1'b1;
        end else begin
            p2_7_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_1_ce0 = 1'b1;
        end else begin
            p2_7_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_7_2_ce0 = 1'b1;
        end else begin
            p2_7_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_0_ce0 = 1'b1;
        end else begin
            p2_8_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_1_ce0 = 1'b1;
        end else begin
            p2_8_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            p2_8_2_ce0 = 1'b1;
        end else begin
            p2_8_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_idle_pp0_1to4 == 1'b1) & (ap_start == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_reset_idle_pp0 == 1'b0))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_reset_idle_pp0 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln120_5_fu_1022_p2 = (sub_ln120_2_fu_1012_p2 + 7'd1);

    assign add_ln120_6_fu_1053_p2 = (sub_ln120_2_reg_3918 + 7'd2);

    assign add_ln120_7_fu_1083_p2 = (mul_ln120_reg_3753 + 7'd1);

    assign add_ln120_8_fu_1163_p2 = (mul_ln120_reg_3753 + 7'd2);

    assign add_ln120_fu_986_p2 = ($signed(
        sext_ln120_fu_982_p1
    ) + $signed(
        axis_offset1_cast3_fu_926_p1
    ));

    assign add_ln129_24_fu_1093_p2 = (mul_ln120_reg_3753 + 7'd4);

    assign add_ln129_25_fu_1173_p2 = (mul_ln120_reg_3753 + 7'd5);

    assign add_ln129_26_fu_1043_p2 = (mul_ln120_reg_3753 + 7'd6);

    assign add_ln129_27_fu_1103_p2 = (mul_ln120_reg_3753 + 7'd7);

    assign add_ln129_28_fu_1203_p2 = (mul_ln120_reg_3753 + 7'd8);

    assign add_ln129_29_fu_1063_p2 = (mul_ln120_reg_3753 + 7'd9);

    assign add_ln129_30_fu_1123_p2 = (mul_ln120_reg_3753 + 7'd10);

    assign add_ln129_31_fu_1223_p2 = (mul_ln120_reg_3753 + 7'd11);

    assign add_ln129_32_fu_1073_p2 = (mul_ln120_reg_3753 + 7'd12);

    assign add_ln129_33_fu_1143_p2 = (mul_ln120_reg_3753 + 7'd13);

    assign add_ln129_34_fu_1243_p2 = (mul_ln120_reg_3753 + 7'd14);

    assign add_ln129_35_fu_1113_p2 = (mul_ln120_reg_3753 + 7'd15);

    assign add_ln129_36_fu_1183_p2 = (mul_ln120_reg_3753 + 7'd16);

    assign add_ln129_37_fu_1263_p2 = (mul_ln120_reg_3753 + 7'd17);

    assign add_ln129_38_fu_1133_p2 = (mul_ln120_reg_3753 + 7'd18);

    assign add_ln129_39_fu_1213_p2 = (mul_ln120_reg_3753 + 7'd19);

    assign add_ln129_40_fu_1273_p2 = (mul_ln120_reg_3753 + 7'd20);

    assign add_ln129_41_fu_1153_p2 = (mul_ln120_reg_3753 + 7'd21);

    assign add_ln129_42_fu_1233_p2 = (mul_ln120_reg_3753 + 7'd22);

    assign add_ln129_43_fu_1283_p2 = (mul_ln120_reg_3753 + 7'd23);

    assign add_ln129_44_fu_1193_p2 = (mul_ln120_reg_3753 + 7'd24);

    assign add_ln129_45_fu_1253_p2 = (mul_ln120_reg_3753 + 7'd25);

    assign add_ln129_46_fu_1293_p2 = (mul_ln120_reg_3753 + 7'd26);

    assign add_ln129_fu_1033_p2 = (mul_ln120_reg_3753 + 7'd3);

    assign and_ln133_16_fu_1381_p2 = (grp_fu_803_p2 & and_ln133_fu_1375_p2);

    assign and_ln133_17_fu_1584_p2 = (or_ln133_18_fu_1578_p2 & or_ln133_17_fu_1560_p2);

    assign and_ln133_18_fu_1590_p2 = (grp_fu_803_p2 & and_ln133_17_fu_1584_p2);

    assign and_ln133_19_fu_1871_p2 = (or_ln133_20_fu_1865_p2 & or_ln133_19_fu_1847_p2);

    assign and_ln133_20_fu_1877_p2 = (grp_fu_803_p2 & and_ln133_19_fu_1871_p2);

    assign and_ln133_21_fu_2158_p2 = (or_ln133_22_fu_2152_p2 & or_ln133_21_fu_2134_p2);

    assign and_ln133_22_fu_2164_p2 = (grp_fu_803_p2 & and_ln133_21_fu_2158_p2);

    assign and_ln133_23_fu_2442_p2 = (or_ln133_24_fu_2436_p2 & or_ln133_23_fu_2418_p2);

    assign and_ln133_24_fu_2448_p2 = (grp_fu_803_p2 & and_ln133_23_fu_2442_p2);

    assign and_ln133_25_fu_2729_p2 = (or_ln133_26_fu_2723_p2 & or_ln133_25_fu_2705_p2);

    assign and_ln133_26_fu_2735_p2 = (grp_fu_803_p2 & and_ln133_25_fu_2729_p2);

    assign and_ln133_27_fu_3016_p2 = (or_ln133_28_fu_3010_p2 & or_ln133_27_fu_2992_p2);

    assign and_ln133_28_fu_3022_p2 = (grp_fu_803_p2 & and_ln133_27_fu_3016_p2);

    assign and_ln133_29_fu_3303_p2 = (or_ln133_30_fu_3297_p2 & or_ln133_29_fu_3279_p2);

    assign and_ln133_30_fu_3309_p2 = (grp_fu_807_p2 & and_ln133_29_fu_3303_p2);

    assign and_ln133_fu_1375_p2 = (or_ln133_fu_1351_p2 & or_ln133_16_fu_1369_p2);

    assign and_ln134_15_fu_1638_p2 = (or_ln134_fu_1632_p2 & or_ln133_17_fu_1560_p2);

    assign and_ln134_16_fu_1644_p2 = (grp_fu_807_p2 & and_ln134_15_fu_1638_p2);

    assign and_ln134_17_fu_1925_p2 = (or_ln134_7_fu_1919_p2 & or_ln133_19_fu_1847_p2);

    assign and_ln134_18_fu_1931_p2 = (grp_fu_807_p2 & and_ln134_17_fu_1925_p2);

    assign and_ln134_19_fu_2212_p2 = (or_ln134_8_fu_2206_p2 & or_ln133_21_fu_2134_p2);

    assign and_ln134_20_fu_2218_p2 = (grp_fu_807_p2 & and_ln134_19_fu_2212_p2);

    assign and_ln134_21_fu_2496_p2 = (or_ln134_9_fu_2490_p2 & or_ln133_23_fu_2418_p2);

    assign and_ln134_22_fu_2502_p2 = (grp_fu_807_p2 & and_ln134_21_fu_2496_p2);

    assign and_ln134_23_fu_2783_p2 = (or_ln134_10_fu_2777_p2 & or_ln133_25_fu_2705_p2);

    assign and_ln134_24_fu_2789_p2 = (grp_fu_807_p2 & and_ln134_23_fu_2783_p2);

    assign and_ln134_25_fu_3070_p2 = (or_ln134_11_fu_3064_p2 & or_ln133_27_fu_2992_p2);

    assign and_ln134_26_fu_3076_p2 = (grp_fu_807_p2 & and_ln134_25_fu_3070_p2);

    assign and_ln134_27_fu_3357_p2 = (or_ln134_12_fu_3351_p2 & or_ln133_29_fu_3279_p2);

    assign and_ln134_28_fu_3363_p2 = (grp_fu_811_p2 & and_ln134_27_fu_3357_p2);

    assign and_ln134_fu_1395_p2 = (grp_fu_807_p2 & and_ln133_fu_1375_p2);

    assign and_ln135_16_fu_1487_p2 = (tmp_93_reg_4742 & and_ln135_reg_4736);

    assign and_ln135_17_fu_1728_p2 = (or_ln135_18_fu_1722_p2 & or_ln135_17_fu_1704_p2);

    assign and_ln135_18_fu_1734_p2 = (grp_fu_811_p2 & and_ln135_17_fu_1728_p2);

    assign and_ln135_19_fu_2015_p2 = (or_ln135_20_fu_2009_p2 & or_ln135_19_fu_1991_p2);

    assign and_ln135_20_fu_2021_p2 = (grp_fu_811_p2 & and_ln135_19_fu_2015_p2);

    assign and_ln135_21_fu_2301_p2 = (or_ln135_22_fu_2295_p2 & or_ln135_21_fu_2277_p2);

    assign and_ln135_22_fu_2307_p2 = (grp_fu_811_p2 & and_ln135_21_fu_2301_p2);

    assign and_ln135_23_fu_2586_p2 = (or_ln135_24_fu_2580_p2 & or_ln135_23_fu_2562_p2);

    assign and_ln135_24_fu_2592_p2 = (grp_fu_811_p2 & and_ln135_23_fu_2586_p2);

    assign and_ln135_25_fu_2873_p2 = (or_ln135_26_fu_2867_p2 & or_ln135_25_fu_2849_p2);

    assign and_ln135_26_fu_2879_p2 = (grp_fu_811_p2 & and_ln135_25_fu_2873_p2);

    assign and_ln135_27_fu_3160_p2 = (or_ln135_28_fu_3154_p2 & or_ln135_27_fu_3136_p2);

    assign and_ln135_28_fu_3166_p2 = (grp_fu_811_p2 & and_ln135_27_fu_3160_p2);

    assign and_ln135_29_fu_3446_p2 = (or_ln135_30_fu_3440_p2 & or_ln135_29_fu_3422_p2);

    assign and_ln135_30_fu_3452_p2 = (grp_fu_807_p2 & and_ln135_29_fu_3446_p2);

    assign and_ln135_fu_1481_p2 = (or_ln135_fu_1457_p2 & or_ln135_16_fu_1475_p2);

    assign and_ln136_15_fu_1782_p2 = (or_ln136_fu_1776_p2 & or_ln135_17_reg_4789);

    assign and_ln136_16_fu_1787_p2 = (grp_fu_803_p2 & and_ln136_15_fu_1782_p2);

    assign and_ln136_17_fu_2069_p2 = (or_ln136_7_fu_2063_p2 & or_ln135_19_reg_4822);

    assign and_ln136_18_fu_2074_p2 = (grp_fu_803_p2 & and_ln136_17_fu_2069_p2);

    assign and_ln136_19_fu_2354_p2 = (or_ln136_8_fu_2348_p2 & or_ln135_21_reg_4855);

    assign and_ln136_20_fu_2359_p2 = (grp_fu_803_p2 & and_ln136_19_fu_2354_p2);

    assign and_ln136_21_fu_2640_p2 = (or_ln136_9_fu_2634_p2 & or_ln135_23_reg_4888);

    assign and_ln136_22_fu_2645_p2 = (grp_fu_803_p2 & and_ln136_21_fu_2640_p2);

    assign and_ln136_23_fu_2927_p2 = (or_ln136_10_fu_2921_p2 & or_ln135_25_reg_4930);

    assign and_ln136_24_fu_2932_p2 = (grp_fu_803_p2 & and_ln136_23_fu_2927_p2);

    assign and_ln136_25_fu_3214_p2 = (or_ln136_11_fu_3208_p2 & or_ln135_27_reg_4963);

    assign and_ln136_26_fu_3219_p2 = (grp_fu_803_p2 & and_ln136_25_fu_3214_p2);

    assign and_ln136_27_fu_3499_p2 = (or_ln136_12_fu_3493_p2 & or_ln135_29_fu_3422_p2);

    assign and_ln136_28_fu_3505_p2 = (grp_fu_811_p2 & and_ln136_27_fu_3499_p2);

    assign and_ln136_fu_1500_p2 = (grp_fu_803_p2 & and_ln135_reg_4736);

    assign and_ln139_5_fu_3587_p2 = (or_ln139_fu_3563_p2 & or_ln139_3_fu_3581_p2);

    assign and_ln139_6_fu_3728_p2 = (tmp_167_reg_5053 & and_ln139_5_reg_5032);

    assign and_ln139_7_fu_3628_p2 = (or_ln139_fu_3563_p2 & or_ln139_4_fu_3622_p2);

    assign and_ln139_8_fu_3634_p2 = (tmp_169_reg_5012 & and_ln139_7_fu_3628_p2);

    assign and_ln139_fu_3732_p2 = (and_ln139_8_reg_5037 & and_ln139_6_fu_3728_p2);

    assign and_ln140_5_fu_3674_p2 = (or_ln140_4_fu_3668_p2 & or_ln139_3_fu_3581_p2);

    assign and_ln140_6_fu_3680_p2 = (tmp_171_reg_5017 & and_ln140_5_fu_3674_p2);

    assign and_ln140_7_fu_3685_p2 = (or_ln140_4_fu_3668_p2 & or_ln139_4_fu_3622_p2);

    assign and_ln140_8_fu_3691_p2 = (tmp_172_reg_5022 & and_ln140_7_fu_3685_p2);

    assign and_ln140_fu_3707_p2 = (or_ln140_fu_3701_p2 & and_ln140_6_fu_3680_p2);

    assign and_ln141_fu_3696_p2 = (tmp_173_reg_5027 & and_ln139_5_fu_3587_p2);

    assign and_ln142_2_fu_3713_p2 = (grp_fu_811_p2 & and_ln140_7_reg_5043);

    assign and_ln142_fu_3718_p2 = (and_ln142_2_fu_3713_p2 & and_ln139_8_reg_5037);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_return = (or_ln140_5_reg_5058 | and_ln139_fu_3732_p2);

    assign axis_address1 = zext_ln120_10_fu_1017_p1;

    assign axis_offset1_cast3_fu_926_p1 = axis_offset1;

    assign bitcast_ln133_16_fu_1321_p1 = reg_886;

    assign bitcast_ln133_17_fu_1513_p1 = reg_901;

    assign bitcast_ln133_18_fu_1531_p1 = max1_reg_4722;

    assign bitcast_ln133_19_fu_1800_p1 = reg_886;

    assign bitcast_ln133_20_fu_1818_p1 = max1_15_reg_4775;

    assign bitcast_ln133_21_fu_2087_p1 = reg_919;

    assign bitcast_ln133_22_fu_2105_p1 = max1_16_reg_4808;

    assign bitcast_ln133_23_fu_2371_p1 = reg_851;

    assign bitcast_ln133_24_fu_2389_p1 = max1_17_reg_4841;

    assign bitcast_ln133_25_fu_2658_p1 = reg_865;

    assign bitcast_ln133_26_fu_2676_p1 = max1_18_reg_4874;

    assign bitcast_ln133_27_fu_2945_p1 = reg_901;

    assign bitcast_ln133_28_fu_2963_p1 = max1_19_reg_4916;

    assign bitcast_ln133_29_fu_3232_p1 = reg_919;

    assign bitcast_ln133_30_fu_3250_p1 = max1_20_reg_4949;

    assign bitcast_ln133_fu_1303_p1 = reg_872;

    assign bitcast_ln134_10_fu_2748_p1 = min1_15_reg_4881;

    assign bitcast_ln134_11_fu_3035_p1 = min1_16_reg_4923;

    assign bitcast_ln134_12_fu_3322_p1 = min1_17_reg_4956;

    assign bitcast_ln134_7_fu_1890_p1 = min1_12_reg_4782;

    assign bitcast_ln134_8_fu_2177_p1 = min1_13_reg_4815;

    assign bitcast_ln134_9_fu_2461_p1 = min1_14_reg_4848;

    assign bitcast_ln134_fu_1603_p1 = min1_11_reg_4729;

    assign bitcast_ln135_16_fu_1427_p1 = reg_894;

    assign bitcast_ln135_17_fu_1657_p1 = reg_907;

    assign bitcast_ln135_18_fu_1675_p1 = max2_reg_4747;

    assign bitcast_ln135_19_fu_1944_p1 = reg_913;

    assign bitcast_ln135_20_fu_1962_p1 = max2_15_reg_4794;

    assign bitcast_ln135_21_fu_2231_p1 = n2_25_reg_4761;

    assign bitcast_ln135_22_fu_2248_p1 = max2_16_reg_4827;

    assign bitcast_ln135_23_fu_2515_p1 = reg_858;

    assign bitcast_ln135_24_fu_2533_p1 = max2_17_reg_4860;

    assign bitcast_ln135_25_fu_2802_p1 = reg_907;

    assign bitcast_ln135_26_fu_2820_p1 = max2_18_reg_4893;

    assign bitcast_ln135_27_fu_3089_p1 = reg_913;

    assign bitcast_ln135_28_fu_3107_p1 = max2_19_reg_4935;

    assign bitcast_ln135_29_fu_3376_p1 = n2_37_reg_4900;

    assign bitcast_ln135_30_fu_3393_p1 = max2_20_reg_4968;

    assign bitcast_ln135_fu_1409_p1 = reg_879;

    assign bitcast_ln136_10_fu_2892_p1 = min2_15_reg_4909;

    assign bitcast_ln136_11_fu_3179_p1 = min2_16_reg_4942;

    assign bitcast_ln136_12_fu_3464_p1 = min2_17_reg_4975;

    assign bitcast_ln136_7_fu_2034_p1 = min2_12_reg_4801;

    assign bitcast_ln136_8_fu_2319_p1 = min2_13_reg_4834;

    assign bitcast_ln136_9_fu_2605_p1 = min2_14_reg_4867;

    assign bitcast_ln136_fu_1747_p1 = min2_11_reg_4754;

    assign bitcast_ln139_3_fu_3534_p1 = max2_21_reg_4997;

    assign bitcast_ln139_4_fu_3593_p1 = min2_18_reg_5005;

    assign bitcast_ln139_fu_3517_p1 = max1_21_reg_4982;

    assign bitcast_ln140_fu_3639_p1 = min1_18_reg_4989;

    assign icmp_ln133_32_fu_1345_p2 = ((trunc_ln133_fu_1317_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_33_fu_1357_p2 = ((tmp_88_fu_1325_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_34_fu_1363_p2 = ((trunc_ln133_16_fu_1335_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_35_fu_1548_p2 = ((tmp_95_fu_1517_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_36_fu_1554_p2 = ((trunc_ln133_17_fu_1527_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_37_fu_1566_p2 = ((tmp_96_fu_1534_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_38_fu_1572_p2 = ((trunc_ln133_18_fu_1544_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_39_fu_1835_p2 = ((tmp_105_fu_1804_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_40_fu_1841_p2 = ((trunc_ln133_19_fu_1814_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_41_fu_1853_p2 = ((tmp_106_fu_1821_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_42_fu_1859_p2 = ((trunc_ln133_20_fu_1831_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_43_fu_2122_p2 = ((tmp_115_fu_2091_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_44_fu_2128_p2 = ((trunc_ln133_21_fu_2101_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_45_fu_2140_p2 = ((tmp_116_fu_2108_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_46_fu_2146_p2 = ((trunc_ln133_22_fu_2118_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_47_fu_2406_p2 = ((tmp_125_fu_2375_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_48_fu_2412_p2 = ((trunc_ln133_23_fu_2385_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_49_fu_2424_p2 = ((tmp_126_fu_2392_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_50_fu_2430_p2 = ((trunc_ln133_24_fu_2402_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_51_fu_2693_p2 = ((tmp_135_fu_2662_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_52_fu_2699_p2 = ((trunc_ln133_25_fu_2672_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_53_fu_2711_p2 = ((tmp_136_fu_2679_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_54_fu_2717_p2 = ((trunc_ln133_26_fu_2689_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_55_fu_2980_p2 = ((tmp_145_fu_2949_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_56_fu_2986_p2 = ((trunc_ln133_27_fu_2959_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_57_fu_2998_p2 = ((tmp_146_fu_2966_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_58_fu_3004_p2 = ((trunc_ln133_28_fu_2976_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_59_fu_3267_p2 = ((tmp_155_fu_3236_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_60_fu_3273_p2 = ((trunc_ln133_29_fu_3246_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_61_fu_3285_p2 = ((tmp_156_fu_3253_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln133_62_fu_3291_p2 = ((trunc_ln133_30_fu_3263_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln133_fu_1339_p2 = ((tmp_s_fu_1307_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_14_fu_1626_p2 = ((trunc_ln134_fu_1616_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_15_fu_1907_p2 = ((tmp_108_fu_1893_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_16_fu_1913_p2 = ((trunc_ln134_7_fu_1903_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_17_fu_2194_p2 = ((tmp_118_fu_2180_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_18_fu_2200_p2 = ((trunc_ln134_8_fu_2190_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_19_fu_2478_p2 = ((tmp_128_fu_2464_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_20_fu_2484_p2 = ((trunc_ln134_9_fu_2474_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_21_fu_2765_p2 = ((tmp_138_fu_2751_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_22_fu_2771_p2 = ((trunc_ln134_10_fu_2761_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_23_fu_3052_p2 = ((tmp_148_fu_3038_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_24_fu_3058_p2 = ((trunc_ln134_11_fu_3048_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_25_fu_3339_p2 = ((tmp_158_fu_3325_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_26_fu_3345_p2 = ((trunc_ln134_12_fu_3335_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln134_fu_1620_p2 = ((tmp_98_fu_1606_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_32_fu_1451_p2 = ((trunc_ln135_fu_1423_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_33_fu_1463_p2 = ((tmp_92_fu_1431_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_34_fu_1469_p2 = ((trunc_ln135_16_fu_1441_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_35_fu_1692_p2 = ((tmp_100_fu_1661_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_36_fu_1698_p2 = ((trunc_ln135_17_fu_1671_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_37_fu_1710_p2 = ((tmp_101_fu_1678_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_38_fu_1716_p2 = ((trunc_ln135_18_fu_1688_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_39_fu_1979_p2 = ((tmp_110_fu_1948_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_40_fu_1985_p2 = ((trunc_ln135_19_fu_1958_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_41_fu_1997_p2 = ((tmp_111_fu_1965_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_42_fu_2003_p2 = ((trunc_ln135_20_fu_1975_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_43_fu_2265_p2 = ((tmp_120_fu_2234_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_44_fu_2271_p2 = ((trunc_ln135_21_fu_2244_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_45_fu_2283_p2 = ((tmp_121_fu_2251_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_46_fu_2289_p2 = ((trunc_ln135_22_fu_2261_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_47_fu_2550_p2 = ((tmp_130_fu_2519_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_48_fu_2556_p2 = ((trunc_ln135_23_fu_2529_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_49_fu_2568_p2 = ((tmp_131_fu_2536_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_50_fu_2574_p2 = ((trunc_ln135_24_fu_2546_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_51_fu_2837_p2 = ((tmp_140_fu_2806_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_52_fu_2843_p2 = ((trunc_ln135_25_fu_2816_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_53_fu_2855_p2 = ((tmp_141_fu_2823_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_54_fu_2861_p2 = ((trunc_ln135_26_fu_2833_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_55_fu_3124_p2 = ((tmp_150_fu_3093_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_56_fu_3130_p2 = ((trunc_ln135_27_fu_3103_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_57_fu_3142_p2 = ((tmp_151_fu_3110_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_58_fu_3148_p2 = ((trunc_ln135_28_fu_3120_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_59_fu_3410_p2 = ((tmp_160_fu_3379_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_60_fu_3416_p2 = ((trunc_ln135_29_fu_3389_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_61_fu_3428_p2 = ((tmp_161_fu_3396_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln135_62_fu_3434_p2 = ((trunc_ln135_30_fu_3406_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln135_fu_1445_p2 = ((tmp_91_fu_1413_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_14_fu_1770_p2 = ((trunc_ln136_fu_1760_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_15_fu_2051_p2 = ((tmp_113_fu_2037_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_16_fu_2057_p2 = ((trunc_ln136_7_fu_2047_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_17_fu_2336_p2 = ((tmp_123_fu_2322_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_18_fu_2342_p2 = ((trunc_ln136_8_fu_2332_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_19_fu_2622_p2 = ((tmp_133_fu_2608_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_20_fu_2628_p2 = ((trunc_ln136_9_fu_2618_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_21_fu_2909_p2 = ((tmp_143_fu_2895_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_22_fu_2915_p2 = ((trunc_ln136_10_fu_2905_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_23_fu_3196_p2 = ((tmp_153_fu_3182_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_24_fu_3202_p2 = ((trunc_ln136_11_fu_3192_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_25_fu_3481_p2 = ((tmp_163_fu_3467_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln136_26_fu_3487_p2 = ((trunc_ln136_12_fu_3477_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln136_fu_1764_p2 = ((tmp_103_fu_1750_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_10_fu_3616_p2 = ((trunc_ln139_4_fu_3606_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_6_fu_3557_p2 = ((trunc_ln139_fu_3530_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_7_fu_3569_p2 = ((tmp_166_fu_3537_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_8_fu_3575_p2 = ((trunc_ln139_3_fu_3547_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln139_9_fu_3610_p2 = ((tmp_168_fu_3596_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln139_fu_3551_p2 = ((tmp_165_fu_3520_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln140_2_fu_3662_p2 = ((trunc_ln140_fu_3652_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln140_fu_3656_p2 = ((tmp_170_fu_3642_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign max1_15_fu_1596_p3 = ((and_ln133_18_fu_1590_p2[0:0] == 1'b1) ? reg_901 : max1_reg_4722);

    assign max1_16_fu_1883_p3 = ((and_ln133_20_fu_1877_p2[0:0] == 1'b1) ? reg_886 : max1_15_reg_4775);

    assign max1_17_fu_2170_p3 = ((and_ln133_22_fu_2164_p2[0:0] == 1'b1) ? reg_919 : max1_16_reg_4808);

    assign max1_18_fu_2454_p3 = ((and_ln133_24_fu_2448_p2[0:0] == 1'b1) ? reg_851 : max1_17_reg_4841);

    assign max1_19_fu_2741_p3 = ((and_ln133_26_fu_2735_p2[0:0] == 1'b1) ? reg_865 : max1_18_reg_4874);

    assign max1_20_fu_3028_p3 = ((and_ln133_28_fu_3022_p2[0:0] == 1'b1) ? reg_901 : max1_19_reg_4916);

    assign max1_21_fu_3315_p3 = ((and_ln133_30_fu_3309_p2[0:0] == 1'b1) ? reg_919 : max1_20_reg_4949);

    assign max1_fu_1387_p3 = ((and_ln133_16_fu_1381_p2[0:0] == 1'b1) ? reg_872 : reg_886);

    assign max2_15_fu_1740_p3 = ((and_ln135_18_fu_1734_p2[0:0] == 1'b1) ? reg_907 : max2_reg_4747);

    assign max2_16_fu_2027_p3 = ((and_ln135_20_fu_2021_p2[0:0] == 1'b1) ? reg_913 : max2_15_reg_4794);

    assign max2_17_fu_2313_p3 = ((and_ln135_22_fu_2307_p2[0:0] == 1'b1) ? n2_25_reg_4761 : max2_16_reg_4827);

    assign max2_18_fu_2598_p3 = ((and_ln135_24_fu_2592_p2[0:0] == 1'b1) ? reg_858 : max2_17_reg_4860);

    assign max2_19_fu_2885_p3 = ((and_ln135_26_fu_2879_p2[0:0] == 1'b1) ? reg_907 : max2_18_reg_4893);

    assign max2_20_fu_3172_p3 = ((and_ln135_28_fu_3166_p2[0:0] == 1'b1) ? reg_913 : max2_19_reg_4935);

    assign max2_21_fu_3458_p3 = ((and_ln135_30_fu_3452_p2[0:0] == 1'b1) ? n2_37_reg_4900 : max2_20_reg_4968);

    assign max2_fu_1491_p3 = ((and_ln135_16_fu_1487_p2[0:0] == 1'b1) ? reg_879 : reg_894);

    assign min1_11_fu_1401_p3 = ((and_ln134_fu_1395_p2[0:0] == 1'b1) ? reg_872 : reg_886);

    assign min1_12_fu_1650_p3 = ((and_ln134_16_fu_1644_p2[0:0] == 1'b1) ? reg_901 : min1_11_reg_4729);

    assign min1_13_fu_1937_p3 = ((and_ln134_18_fu_1931_p2[0:0] == 1'b1) ? reg_886 : min1_12_reg_4782);

    assign min1_14_fu_2224_p3 = ((and_ln134_20_fu_2218_p2[0:0] == 1'b1) ? reg_919 : min1_13_reg_4815);

    assign min1_15_fu_2508_p3 = ((and_ln134_22_fu_2502_p2[0:0] == 1'b1) ? reg_851 : min1_14_reg_4848);

    assign min1_16_fu_2795_p3 = ((and_ln134_24_fu_2789_p2[0:0] == 1'b1) ? reg_865 : min1_15_reg_4881);

    assign min1_17_fu_3082_p3 = ((and_ln134_26_fu_3076_p2[0:0] == 1'b1) ? reg_901 : min1_16_reg_4923);

    assign min1_18_fu_3369_p3 = ((and_ln134_28_fu_3363_p2[0:0] == 1'b1) ? reg_919 : min1_17_reg_4956);

    assign min2_11_fu_1505_p3 = ((and_ln136_fu_1500_p2[0:0] == 1'b1) ? reg_879 : reg_894);

    assign min2_12_fu_1793_p3 = ((and_ln136_16_fu_1787_p2[0:0] == 1'b1) ? reg_907 : min2_11_reg_4754);

    assign min2_13_fu_2080_p3 = ((and_ln136_18_fu_2074_p2[0:0] == 1'b1) ? reg_913 : min2_12_reg_4801);

    assign min2_14_fu_2365_p3 = ((and_ln136_20_fu_2359_p2[0:0] == 1'b1) ? n2_25_reg_4761 : min2_13_reg_4834);

    assign min2_15_fu_2651_p3 = ((and_ln136_22_fu_2645_p2[0:0] == 1'b1) ? reg_858 : min2_14_reg_4867);

    assign min2_16_fu_2938_p3 = ((and_ln136_24_fu_2932_p2[0:0] == 1'b1) ? reg_907 : min2_15_reg_4909);

    assign min2_17_fu_3225_p3 = ((and_ln136_26_fu_3219_p2[0:0] == 1'b1) ? reg_913 : min2_16_reg_4942);

    assign min2_18_fu_3511_p3 = ((and_ln136_28_fu_3505_p2[0:0] == 1'b1) ? n2_37_reg_4900 : min2_17_reg_4975);

    assign mul_ln120_fu_996_p0 = mul_ln120_fu_996_p00;

    assign mul_ln120_fu_996_p00 = p1_offset;

    assign mul_ln120_fu_996_p1 = 7'd27;

    assign or_ln133_16_fu_1369_p2 = (icmp_ln133_34_fu_1363_p2 | icmp_ln133_33_fu_1357_p2);

    assign or_ln133_17_fu_1560_p2 = (icmp_ln133_36_fu_1554_p2 | icmp_ln133_35_fu_1548_p2);

    assign or_ln133_18_fu_1578_p2 = (icmp_ln133_38_fu_1572_p2 | icmp_ln133_37_fu_1566_p2);

    assign or_ln133_19_fu_1847_p2 = (icmp_ln133_40_fu_1841_p2 | icmp_ln133_39_fu_1835_p2);

    assign or_ln133_20_fu_1865_p2 = (icmp_ln133_42_fu_1859_p2 | icmp_ln133_41_fu_1853_p2);

    assign or_ln133_21_fu_2134_p2 = (icmp_ln133_44_fu_2128_p2 | icmp_ln133_43_fu_2122_p2);

    assign or_ln133_22_fu_2152_p2 = (icmp_ln133_46_fu_2146_p2 | icmp_ln133_45_fu_2140_p2);

    assign or_ln133_23_fu_2418_p2 = (icmp_ln133_48_fu_2412_p2 | icmp_ln133_47_fu_2406_p2);

    assign or_ln133_24_fu_2436_p2 = (icmp_ln133_50_fu_2430_p2 | icmp_ln133_49_fu_2424_p2);

    assign or_ln133_25_fu_2705_p2 = (icmp_ln133_52_fu_2699_p2 | icmp_ln133_51_fu_2693_p2);

    assign or_ln133_26_fu_2723_p2 = (icmp_ln133_54_fu_2717_p2 | icmp_ln133_53_fu_2711_p2);

    assign or_ln133_27_fu_2992_p2 = (icmp_ln133_56_fu_2986_p2 | icmp_ln133_55_fu_2980_p2);

    assign or_ln133_28_fu_3010_p2 = (icmp_ln133_58_fu_3004_p2 | icmp_ln133_57_fu_2998_p2);

    assign or_ln133_29_fu_3279_p2 = (icmp_ln133_60_fu_3273_p2 | icmp_ln133_59_fu_3267_p2);

    assign or_ln133_30_fu_3297_p2 = (icmp_ln133_62_fu_3291_p2 | icmp_ln133_61_fu_3285_p2);

    assign or_ln133_fu_1351_p2 = (icmp_ln133_fu_1339_p2 | icmp_ln133_32_fu_1345_p2);

    assign or_ln134_10_fu_2777_p2 = (icmp_ln134_22_fu_2771_p2 | icmp_ln134_21_fu_2765_p2);

    assign or_ln134_11_fu_3064_p2 = (icmp_ln134_24_fu_3058_p2 | icmp_ln134_23_fu_3052_p2);

    assign or_ln134_12_fu_3351_p2 = (icmp_ln134_26_fu_3345_p2 | icmp_ln134_25_fu_3339_p2);

    assign or_ln134_7_fu_1919_p2 = (icmp_ln134_16_fu_1913_p2 | icmp_ln134_15_fu_1907_p2);

    assign or_ln134_8_fu_2206_p2 = (icmp_ln134_18_fu_2200_p2 | icmp_ln134_17_fu_2194_p2);

    assign or_ln134_9_fu_2490_p2 = (icmp_ln134_20_fu_2484_p2 | icmp_ln134_19_fu_2478_p2);

    assign or_ln134_fu_1632_p2 = (icmp_ln134_fu_1620_p2 | icmp_ln134_14_fu_1626_p2);

    assign or_ln135_16_fu_1475_p2 = (icmp_ln135_34_fu_1469_p2 | icmp_ln135_33_fu_1463_p2);

    assign or_ln135_17_fu_1704_p2 = (icmp_ln135_36_fu_1698_p2 | icmp_ln135_35_fu_1692_p2);

    assign or_ln135_18_fu_1722_p2 = (icmp_ln135_38_fu_1716_p2 | icmp_ln135_37_fu_1710_p2);

    assign or_ln135_19_fu_1991_p2 = (icmp_ln135_40_fu_1985_p2 | icmp_ln135_39_fu_1979_p2);

    assign or_ln135_20_fu_2009_p2 = (icmp_ln135_42_fu_2003_p2 | icmp_ln135_41_fu_1997_p2);

    assign or_ln135_21_fu_2277_p2 = (icmp_ln135_44_fu_2271_p2 | icmp_ln135_43_fu_2265_p2);

    assign or_ln135_22_fu_2295_p2 = (icmp_ln135_46_fu_2289_p2 | icmp_ln135_45_fu_2283_p2);

    assign or_ln135_23_fu_2562_p2 = (icmp_ln135_48_fu_2556_p2 | icmp_ln135_47_fu_2550_p2);

    assign or_ln135_24_fu_2580_p2 = (icmp_ln135_50_fu_2574_p2 | icmp_ln135_49_fu_2568_p2);

    assign or_ln135_25_fu_2849_p2 = (icmp_ln135_52_fu_2843_p2 | icmp_ln135_51_fu_2837_p2);

    assign or_ln135_26_fu_2867_p2 = (icmp_ln135_54_fu_2861_p2 | icmp_ln135_53_fu_2855_p2);

    assign or_ln135_27_fu_3136_p2 = (icmp_ln135_56_fu_3130_p2 | icmp_ln135_55_fu_3124_p2);

    assign or_ln135_28_fu_3154_p2 = (icmp_ln135_58_fu_3148_p2 | icmp_ln135_57_fu_3142_p2);

    assign or_ln135_29_fu_3422_p2 = (icmp_ln135_60_fu_3416_p2 | icmp_ln135_59_fu_3410_p2);

    assign or_ln135_30_fu_3440_p2 = (icmp_ln135_62_fu_3434_p2 | icmp_ln135_61_fu_3428_p2);

    assign or_ln135_fu_1457_p2 = (icmp_ln135_fu_1445_p2 | icmp_ln135_32_fu_1451_p2);

    assign or_ln136_10_fu_2921_p2 = (icmp_ln136_22_fu_2915_p2 | icmp_ln136_21_fu_2909_p2);

    assign or_ln136_11_fu_3208_p2 = (icmp_ln136_24_fu_3202_p2 | icmp_ln136_23_fu_3196_p2);

    assign or_ln136_12_fu_3493_p2 = (icmp_ln136_26_fu_3487_p2 | icmp_ln136_25_fu_3481_p2);

    assign or_ln136_7_fu_2063_p2 = (icmp_ln136_16_fu_2057_p2 | icmp_ln136_15_fu_2051_p2);

    assign or_ln136_8_fu_2348_p2 = (icmp_ln136_18_fu_2342_p2 | icmp_ln136_17_fu_2336_p2);

    assign or_ln136_9_fu_2634_p2 = (icmp_ln136_20_fu_2628_p2 | icmp_ln136_19_fu_2622_p2);

    assign or_ln136_fu_1776_p2 = (icmp_ln136_fu_1764_p2 | icmp_ln136_14_fu_1770_p2);

    assign or_ln139_3_fu_3581_p2 = (icmp_ln139_8_fu_3575_p2 | icmp_ln139_7_fu_3569_p2);

    assign or_ln139_4_fu_3622_p2 = (icmp_ln139_9_fu_3610_p2 | icmp_ln139_10_fu_3616_p2);

    assign or_ln139_fu_3563_p2 = (icmp_ln139_fu_3551_p2 | icmp_ln139_6_fu_3557_p2);

    assign or_ln140_4_fu_3668_p2 = (icmp_ln140_fu_3656_p2 | icmp_ln140_2_fu_3662_p2);

    assign or_ln140_5_fu_3723_p2 = (and_ln142_fu_3718_p2 | and_ln140_reg_5048);

    assign or_ln140_fu_3701_p2 = (and_ln141_fu_3696_p2 | and_ln140_8_fu_3691_p2);

    assign p2_0_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_0_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_0_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_1_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_1_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_1_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_2_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_2_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_2_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_3_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_3_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_3_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_4_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_4_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_4_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_5_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_5_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_5_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_6_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_6_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_6_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_7_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_7_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_7_2_address0 = p2_offset_cast_fu_930_p1;

    assign p2_8_0_address0 = p2_offset_cast_fu_930_p1;

    assign p2_8_1_address0 = p2_offset_cast_fu_930_p1;

    assign p2_8_2_address0 = p2_offset_cast_reg_3742;

    assign p2_offset_cast_fu_930_p1 = p2_offset;

    assign sext_ln120_fu_982_p1 = $signed(sub_ln120_fu_976_p2);

    assign shl_ln120_fu_1007_p2 = add_ln120_reg_3747 << 7'd2;

    assign sub_ln120_2_fu_1012_p2 = (shl_ln120_fu_1007_p2 - add_ln120_reg_3747);

    assign sub_ln120_fu_976_p2 = (zext_ln120_9_fu_972_p1 - zext_ln120_fu_960_p1);

    assign tmp_100_fu_1661_p4 = {{bitcast_ln135_17_fu_1657_p1[62:52]}};

    assign tmp_101_fu_1678_p4 = {{bitcast_ln135_18_fu_1675_p1[62:52]}};

    assign tmp_103_fu_1750_p4 = {{bitcast_ln136_fu_1747_p1[62:52]}};

    assign tmp_105_fu_1804_p4 = {{bitcast_ln133_19_fu_1800_p1[62:52]}};

    assign tmp_106_fu_1821_p4 = {{bitcast_ln133_20_fu_1818_p1[62:52]}};

    assign tmp_108_fu_1893_p4 = {{bitcast_ln134_7_fu_1890_p1[62:52]}};

    assign tmp_110_fu_1948_p4 = {{bitcast_ln135_19_fu_1944_p1[62:52]}};

    assign tmp_111_fu_1965_p4 = {{bitcast_ln135_20_fu_1962_p1[62:52]}};

    assign tmp_113_fu_2037_p4 = {{bitcast_ln136_7_fu_2034_p1[62:52]}};

    assign tmp_115_fu_2091_p4 = {{bitcast_ln133_21_fu_2087_p1[62:52]}};

    assign tmp_116_fu_2108_p4 = {{bitcast_ln133_22_fu_2105_p1[62:52]}};

    assign tmp_118_fu_2180_p4 = {{bitcast_ln134_8_fu_2177_p1[62:52]}};

    assign tmp_120_fu_2234_p4 = {{bitcast_ln135_21_fu_2231_p1[62:52]}};

    assign tmp_121_fu_2251_p4 = {{bitcast_ln135_22_fu_2248_p1[62:52]}};

    assign tmp_123_fu_2322_p4 = {{bitcast_ln136_8_fu_2319_p1[62:52]}};

    assign tmp_125_fu_2375_p4 = {{bitcast_ln133_23_fu_2371_p1[62:52]}};

    assign tmp_126_fu_2392_p4 = {{bitcast_ln133_24_fu_2389_p1[62:52]}};

    assign tmp_128_fu_2464_p4 = {{bitcast_ln134_9_fu_2461_p1[62:52]}};

    assign tmp_130_fu_2519_p4 = {{bitcast_ln135_23_fu_2515_p1[62:52]}};

    assign tmp_131_fu_2536_p4 = {{bitcast_ln135_24_fu_2533_p1[62:52]}};

    assign tmp_133_fu_2608_p4 = {{bitcast_ln136_9_fu_2605_p1[62:52]}};

    assign tmp_135_fu_2662_p4 = {{bitcast_ln133_25_fu_2658_p1[62:52]}};

    assign tmp_136_fu_2679_p4 = {{bitcast_ln133_26_fu_2676_p1[62:52]}};

    assign tmp_138_fu_2751_p4 = {{bitcast_ln134_10_fu_2748_p1[62:52]}};

    assign tmp_140_fu_2806_p4 = {{bitcast_ln135_25_fu_2802_p1[62:52]}};

    assign tmp_141_fu_2823_p4 = {{bitcast_ln135_26_fu_2820_p1[62:52]}};

    assign tmp_143_fu_2895_p4 = {{bitcast_ln136_10_fu_2892_p1[62:52]}};

    assign tmp_145_fu_2949_p4 = {{bitcast_ln133_27_fu_2945_p1[62:52]}};

    assign tmp_146_fu_2966_p4 = {{bitcast_ln133_28_fu_2963_p1[62:52]}};

    assign tmp_148_fu_3038_p4 = {{bitcast_ln134_11_fu_3035_p1[62:52]}};

    assign tmp_150_fu_3093_p4 = {{bitcast_ln135_27_fu_3089_p1[62:52]}};

    assign tmp_151_fu_3110_p4 = {{bitcast_ln135_28_fu_3107_p1[62:52]}};

    assign tmp_153_fu_3182_p4 = {{bitcast_ln136_11_fu_3179_p1[62:52]}};

    assign tmp_155_fu_3236_p4 = {{bitcast_ln133_29_fu_3232_p1[62:52]}};

    assign tmp_156_fu_3253_p4 = {{bitcast_ln133_30_fu_3250_p1[62:52]}};

    assign tmp_158_fu_3325_p4 = {{bitcast_ln134_12_fu_3322_p1[62:52]}};

    assign tmp_160_fu_3379_p4 = {{bitcast_ln135_29_fu_3376_p1[62:52]}};

    assign tmp_161_fu_3396_p4 = {{bitcast_ln135_30_fu_3393_p1[62:52]}};

    assign tmp_163_fu_3467_p4 = {{bitcast_ln136_12_fu_3464_p1[62:52]}};

    assign tmp_165_fu_3520_p4 = {{bitcast_ln139_fu_3517_p1[62:52]}};

    assign tmp_166_fu_3537_p4 = {{bitcast_ln139_3_fu_3534_p1[62:52]}};

    assign tmp_168_fu_3596_p4 = {{bitcast_ln139_4_fu_3593_p1[62:52]}};

    assign tmp_170_fu_3642_p4 = {{bitcast_ln140_fu_3639_p1[62:52]}};

    assign tmp_88_fu_1325_p4 = {{bitcast_ln133_16_fu_1321_p1[62:52]}};

    assign tmp_91_fu_1413_p4 = {{bitcast_ln135_fu_1409_p1[62:52]}};

    assign tmp_92_fu_1431_p4 = {{bitcast_ln135_16_fu_1427_p1[62:52]}};

    assign tmp_95_fu_1517_p4 = {{bitcast_ln133_17_fu_1513_p1[62:52]}};

    assign tmp_96_fu_1534_p4 = {{bitcast_ln133_18_fu_1531_p1[62:52]}};

    assign tmp_98_fu_1606_p4 = {{bitcast_ln134_fu_1603_p1[62:52]}};

    assign tmp_fu_964_p3 = {{p2_offset}, {2'd0}};

    assign tmp_s_fu_1307_p4 = {{bitcast_ln133_fu_1303_p1[62:52]}};

    assign trunc_ln133_16_fu_1335_p1 = bitcast_ln133_16_fu_1321_p1[51:0];

    assign trunc_ln133_17_fu_1527_p1 = bitcast_ln133_17_fu_1513_p1[51:0];

    assign trunc_ln133_18_fu_1544_p1 = bitcast_ln133_18_fu_1531_p1[51:0];

    assign trunc_ln133_19_fu_1814_p1 = bitcast_ln133_19_fu_1800_p1[51:0];

    assign trunc_ln133_20_fu_1831_p1 = bitcast_ln133_20_fu_1818_p1[51:0];

    assign trunc_ln133_21_fu_2101_p1 = bitcast_ln133_21_fu_2087_p1[51:0];

    assign trunc_ln133_22_fu_2118_p1 = bitcast_ln133_22_fu_2105_p1[51:0];

    assign trunc_ln133_23_fu_2385_p1 = bitcast_ln133_23_fu_2371_p1[51:0];

    assign trunc_ln133_24_fu_2402_p1 = bitcast_ln133_24_fu_2389_p1[51:0];

    assign trunc_ln133_25_fu_2672_p1 = bitcast_ln133_25_fu_2658_p1[51:0];

    assign trunc_ln133_26_fu_2689_p1 = bitcast_ln133_26_fu_2676_p1[51:0];

    assign trunc_ln133_27_fu_2959_p1 = bitcast_ln133_27_fu_2945_p1[51:0];

    assign trunc_ln133_28_fu_2976_p1 = bitcast_ln133_28_fu_2963_p1[51:0];

    assign trunc_ln133_29_fu_3246_p1 = bitcast_ln133_29_fu_3232_p1[51:0];

    assign trunc_ln133_30_fu_3263_p1 = bitcast_ln133_30_fu_3250_p1[51:0];

    assign trunc_ln133_fu_1317_p1 = bitcast_ln133_fu_1303_p1[51:0];

    assign trunc_ln134_10_fu_2761_p1 = bitcast_ln134_10_fu_2748_p1[51:0];

    assign trunc_ln134_11_fu_3048_p1 = bitcast_ln134_11_fu_3035_p1[51:0];

    assign trunc_ln134_12_fu_3335_p1 = bitcast_ln134_12_fu_3322_p1[51:0];

    assign trunc_ln134_7_fu_1903_p1 = bitcast_ln134_7_fu_1890_p1[51:0];

    assign trunc_ln134_8_fu_2190_p1 = bitcast_ln134_8_fu_2177_p1[51:0];

    assign trunc_ln134_9_fu_2474_p1 = bitcast_ln134_9_fu_2461_p1[51:0];

    assign trunc_ln134_fu_1616_p1 = bitcast_ln134_fu_1603_p1[51:0];

    assign trunc_ln135_16_fu_1441_p1 = bitcast_ln135_16_fu_1427_p1[51:0];

    assign trunc_ln135_17_fu_1671_p1 = bitcast_ln135_17_fu_1657_p1[51:0];

    assign trunc_ln135_18_fu_1688_p1 = bitcast_ln135_18_fu_1675_p1[51:0];

    assign trunc_ln135_19_fu_1958_p1 = bitcast_ln135_19_fu_1944_p1[51:0];

    assign trunc_ln135_20_fu_1975_p1 = bitcast_ln135_20_fu_1962_p1[51:0];

    assign trunc_ln135_21_fu_2244_p1 = bitcast_ln135_21_fu_2231_p1[51:0];

    assign trunc_ln135_22_fu_2261_p1 = bitcast_ln135_22_fu_2248_p1[51:0];

    assign trunc_ln135_23_fu_2529_p1 = bitcast_ln135_23_fu_2515_p1[51:0];

    assign trunc_ln135_24_fu_2546_p1 = bitcast_ln135_24_fu_2533_p1[51:0];

    assign trunc_ln135_25_fu_2816_p1 = bitcast_ln135_25_fu_2802_p1[51:0];

    assign trunc_ln135_26_fu_2833_p1 = bitcast_ln135_26_fu_2820_p1[51:0];

    assign trunc_ln135_27_fu_3103_p1 = bitcast_ln135_27_fu_3089_p1[51:0];

    assign trunc_ln135_28_fu_3120_p1 = bitcast_ln135_28_fu_3107_p1[51:0];

    assign trunc_ln135_29_fu_3389_p1 = bitcast_ln135_29_fu_3376_p1[51:0];

    assign trunc_ln135_30_fu_3406_p1 = bitcast_ln135_30_fu_3393_p1[51:0];

    assign trunc_ln135_fu_1423_p1 = bitcast_ln135_fu_1409_p1[51:0];

    assign trunc_ln136_10_fu_2905_p1 = bitcast_ln136_10_fu_2892_p1[51:0];

    assign trunc_ln136_11_fu_3192_p1 = bitcast_ln136_11_fu_3179_p1[51:0];

    assign trunc_ln136_12_fu_3477_p1 = bitcast_ln136_12_fu_3464_p1[51:0];

    assign trunc_ln136_7_fu_2047_p1 = bitcast_ln136_7_fu_2034_p1[51:0];

    assign trunc_ln136_8_fu_2332_p1 = bitcast_ln136_8_fu_2319_p1[51:0];

    assign trunc_ln136_9_fu_2618_p1 = bitcast_ln136_9_fu_2605_p1[51:0];

    assign trunc_ln136_fu_1760_p1 = bitcast_ln136_fu_1747_p1[51:0];

    assign trunc_ln139_3_fu_3547_p1 = bitcast_ln139_3_fu_3534_p1[51:0];

    assign trunc_ln139_4_fu_3606_p1 = bitcast_ln139_4_fu_3593_p1[51:0];

    assign trunc_ln139_fu_3530_p1 = bitcast_ln139_fu_3517_p1[51:0];

    assign trunc_ln140_fu_3652_p1 = bitcast_ln140_fu_3639_p1[51:0];

    assign zext_ln120_10_fu_1017_p1 = sub_ln120_2_fu_1012_p2;

    assign zext_ln120_11_fu_1028_p1 = add_ln120_5_fu_1022_p2;

    assign zext_ln120_12_fu_1058_p1 = add_ln120_6_fu_1053_p2;

    assign zext_ln120_14_fu_1002_p1 = mul_ln120_fu_996_p2;

    assign zext_ln120_15_fu_1088_p1 = add_ln120_7_fu_1083_p2;

    assign zext_ln120_16_fu_1168_p1 = add_ln120_8_fu_1163_p2;

    assign zext_ln120_9_fu_972_p1 = tmp_fu_964_p3;

    assign zext_ln120_fu_960_p1 = p2_offset;

    assign zext_ln129_24_fu_1098_p1 = add_ln129_24_fu_1093_p2;

    assign zext_ln129_25_fu_1178_p1 = add_ln129_25_fu_1173_p2;

    assign zext_ln129_26_fu_1048_p1 = add_ln129_26_fu_1043_p2;

    assign zext_ln129_27_fu_1108_p1 = add_ln129_27_fu_1103_p2;

    assign zext_ln129_28_fu_1208_p1 = add_ln129_28_fu_1203_p2;

    assign zext_ln129_29_fu_1068_p1 = add_ln129_29_fu_1063_p2;

    assign zext_ln129_30_fu_1128_p1 = add_ln129_30_fu_1123_p2;

    assign zext_ln129_31_fu_1228_p1 = add_ln129_31_fu_1223_p2;

    assign zext_ln129_32_fu_1078_p1 = add_ln129_32_fu_1073_p2;

    assign zext_ln129_33_fu_1148_p1 = add_ln129_33_fu_1143_p2;

    assign zext_ln129_34_fu_1248_p1 = add_ln129_34_fu_1243_p2;

    assign zext_ln129_35_fu_1118_p1 = add_ln129_35_fu_1113_p2;

    assign zext_ln129_36_fu_1188_p1 = add_ln129_36_fu_1183_p2;

    assign zext_ln129_37_fu_1268_p1 = add_ln129_37_fu_1263_p2;

    assign zext_ln129_38_fu_1138_p1 = add_ln129_38_fu_1133_p2;

    assign zext_ln129_39_fu_1218_p1 = add_ln129_39_fu_1213_p2;

    assign zext_ln129_40_fu_1278_p1 = add_ln129_40_fu_1273_p2;

    assign zext_ln129_41_fu_1158_p1 = add_ln129_41_fu_1153_p2;

    assign zext_ln129_42_fu_1238_p1 = add_ln129_42_fu_1233_p2;

    assign zext_ln129_43_fu_1288_p1 = add_ln129_43_fu_1283_p2;

    assign zext_ln129_44_fu_1198_p1 = add_ln129_44_fu_1193_p2;

    assign zext_ln129_45_fu_1258_p1 = add_ln129_45_fu_1253_p2;

    assign zext_ln129_46_fu_1298_p1 = add_ln129_46_fu_1293_p2;

    assign zext_ln129_fu_1038_p1 = add_ln129_fu_1033_p2;

    always @(posedge ap_clk) begin
        p2_offset_cast_reg_3742[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_pointsOverlap_double_1
