/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_57_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    tmp_3,
    empty,
    measurement,
    dx,
    dy,
    ogm_grid_address0,
    ogm_grid_ce0,
    ogm_grid_we0,
    ogm_grid_d0,
    ogm_grid_q0,
    grp_fu_172_p_din0,
    grp_fu_172_p_din1,
    grp_fu_172_p_opcode,
    grp_fu_172_p_dout0,
    grp_fu_172_p_ce,
    grp_fu_194_p_din0,
    grp_fu_194_p_din1,
    grp_fu_194_p_dout0,
    grp_fu_194_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 69'd1;
    parameter ap_ST_fsm_pp0_stage1 = 69'd2;
    parameter ap_ST_fsm_pp0_stage2 = 69'd4;
    parameter ap_ST_fsm_pp0_stage3 = 69'd8;
    parameter ap_ST_fsm_pp0_stage4 = 69'd16;
    parameter ap_ST_fsm_pp0_stage5 = 69'd32;
    parameter ap_ST_fsm_pp0_stage6 = 69'd64;
    parameter ap_ST_fsm_pp0_stage7 = 69'd128;
    parameter ap_ST_fsm_pp0_stage8 = 69'd256;
    parameter ap_ST_fsm_pp0_stage9 = 69'd512;
    parameter ap_ST_fsm_pp0_stage10 = 69'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 69'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 69'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 69'd8192;
    parameter ap_ST_fsm_pp0_stage14 = 69'd16384;
    parameter ap_ST_fsm_pp0_stage15 = 69'd32768;
    parameter ap_ST_fsm_pp0_stage16 = 69'd65536;
    parameter ap_ST_fsm_pp0_stage17 = 69'd131072;
    parameter ap_ST_fsm_pp0_stage18 = 69'd262144;
    parameter ap_ST_fsm_pp0_stage19 = 69'd524288;
    parameter ap_ST_fsm_pp0_stage20 = 69'd1048576;
    parameter ap_ST_fsm_pp0_stage21 = 69'd2097152;
    parameter ap_ST_fsm_pp0_stage22 = 69'd4194304;
    parameter ap_ST_fsm_pp0_stage23 = 69'd8388608;
    parameter ap_ST_fsm_pp0_stage24 = 69'd16777216;
    parameter ap_ST_fsm_pp0_stage25 = 69'd33554432;
    parameter ap_ST_fsm_pp0_stage26 = 69'd67108864;
    parameter ap_ST_fsm_pp0_stage27 = 69'd134217728;
    parameter ap_ST_fsm_pp0_stage28 = 69'd268435456;
    parameter ap_ST_fsm_pp0_stage29 = 69'd536870912;
    parameter ap_ST_fsm_pp0_stage30 = 69'd1073741824;
    parameter ap_ST_fsm_pp0_stage31 = 69'd2147483648;
    parameter ap_ST_fsm_pp0_stage32 = 69'd4294967296;
    parameter ap_ST_fsm_pp0_stage33 = 69'd8589934592;
    parameter ap_ST_fsm_pp0_stage34 = 69'd17179869184;
    parameter ap_ST_fsm_pp0_stage35 = 69'd34359738368;
    parameter ap_ST_fsm_pp0_stage36 = 69'd68719476736;
    parameter ap_ST_fsm_pp0_stage37 = 69'd137438953472;
    parameter ap_ST_fsm_pp0_stage38 = 69'd274877906944;
    parameter ap_ST_fsm_pp0_stage39 = 69'd549755813888;
    parameter ap_ST_fsm_pp0_stage40 = 69'd1099511627776;
    parameter ap_ST_fsm_pp0_stage41 = 69'd2199023255552;
    parameter ap_ST_fsm_pp0_stage42 = 69'd4398046511104;
    parameter ap_ST_fsm_pp0_stage43 = 69'd8796093022208;
    parameter ap_ST_fsm_pp0_stage44 = 69'd17592186044416;
    parameter ap_ST_fsm_pp0_stage45 = 69'd35184372088832;
    parameter ap_ST_fsm_pp0_stage46 = 69'd70368744177664;
    parameter ap_ST_fsm_pp0_stage47 = 69'd140737488355328;
    parameter ap_ST_fsm_pp0_stage48 = 69'd281474976710656;
    parameter ap_ST_fsm_pp0_stage49 = 69'd562949953421312;
    parameter ap_ST_fsm_pp0_stage50 = 69'd1125899906842624;
    parameter ap_ST_fsm_pp0_stage51 = 69'd2251799813685248;
    parameter ap_ST_fsm_pp0_stage52 = 69'd4503599627370496;
    parameter ap_ST_fsm_pp0_stage53 = 69'd9007199254740992;
    parameter ap_ST_fsm_pp0_stage54 = 69'd18014398509481984;
    parameter ap_ST_fsm_pp0_stage55 = 69'd36028797018963968;
    parameter ap_ST_fsm_pp0_stage56 = 69'd72057594037927936;
    parameter ap_ST_fsm_pp0_stage57 = 69'd144115188075855872;
    parameter ap_ST_fsm_pp0_stage58 = 69'd288230376151711744;
    parameter ap_ST_fsm_pp0_stage59 = 69'd576460752303423488;
    parameter ap_ST_fsm_pp0_stage60 = 69'd1152921504606846976;
    parameter ap_ST_fsm_pp0_stage61 = 69'd2305843009213693952;
    parameter ap_ST_fsm_pp0_stage62 = 69'd4611686018427387904;
    parameter ap_ST_fsm_pp0_stage63 = 69'd9223372036854775808;
    parameter ap_ST_fsm_pp0_stage64 = 69'd18446744073709551616;
    parameter ap_ST_fsm_pp0_stage65 = 69'd36893488147419103232;
    parameter ap_ST_fsm_pp0_stage66 = 69'd73786976294838206464;
    parameter ap_ST_fsm_pp0_stage67 = 69'd147573952589676412928;
    parameter ap_ST_fsm_pp0_stage68 = 69'd295147905179352825856;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [10:0] tmp_3;
    input [51:0] empty;
    input [63:0] measurement;
    input [63:0] dx;
    input [63:0] dy;
    output [13:0] ogm_grid_address0;
    output ogm_grid_ce0;
    output ogm_grid_we0;
    output [63:0] ogm_grid_d0;
    input [63:0] ogm_grid_q0;
    output [63:0] grp_fu_172_p_din0;
    output [63:0] grp_fu_172_p_din1;
    output [1:0] grp_fu_172_p_opcode;
    input [63:0] grp_fu_172_p_dout0;
    output grp_fu_172_p_ce;
    output [63:0] grp_fu_194_p_din0;
    output [63:0] grp_fu_194_p_din1;
    input [63:0] grp_fu_194_p_dout0;
    output grp_fu_194_p_ce;

    reg ap_idle;
    reg[13:0] ogm_grid_address0;
    reg ogm_grid_ce0;
    reg ogm_grid_we0;

    (* fsm_encoding = "none" *) reg   [68:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage27;
    wire    ap_block_pp0_stage27_subdone;
    reg   [0:0] and_ln57_1_reg_600;
    reg    ap_condition_exit_pp0_iter0_stage27;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_CS_fsm_pp0_stage68;
    wire    ap_block_pp0_stage68_subdone;
    reg   [63:0] reg_151;
    wire    ap_CS_fsm_pp0_stage20;
    wire    ap_block_pp0_stage20_11001;
    wire    ap_CS_fsm_pp0_stage21;
    wire    ap_block_pp0_stage21_11001;
    wire    ap_block_pp0_stage0_11001;
    wire   [0:0] icmp_ln57_2_fu_164_p2;
    reg   [0:0] icmp_ln57_2_reg_578;
    wire   [0:0] icmp_ln57_3_fu_170_p2;
    reg   [0:0] icmp_ln57_3_reg_583;
    wire   [31:0] i_5_fu_176_p2;
    reg   [31:0] i_5_reg_588;
    wire   [63:0] grp_fu_148_p1;
    reg   [63:0] conv_i_reg_593;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire   [0:0] and_ln57_1_fu_227_p2;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire   [63:0] grp_fu_135_p2;
    reg   [63:0] mul_i_reg_604;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_11001;
    reg   [63:0] mul5_i_reg_609;
    wire    ap_CS_fsm_pp0_stage14;
    wire    ap_block_pp0_stage14_11001;
    reg   [0:0] xs_sign_reg_614;
    wire   [136:0] zext_ln15_fu_273_p1;
    reg   [136:0] zext_ln15_reg_619;
    wire   [0:0] tmp_20_fu_287_p3;
    reg   [0:0] tmp_20_reg_624;
    wire   [136:0] zext_ln18_fu_317_p1;
    reg   [136:0] zext_ln18_reg_629;
    reg   [31:0] tmp_s_reg_634;
    wire   [31:0] val_fu_351_p3;
    reg   [31:0] val_reg_639;
    wire    ap_CS_fsm_pp0_stage22;
    wire    ap_block_pp0_stage22_11001;
    wire   [31:0] result_fu_362_p3;
    reg   [31:0] result_reg_645;
    wire    ap_CS_fsm_pp0_stage23;
    wire    ap_block_pp0_stage23_11001;
    reg   [0:0] xs_sign_1_reg_651;
    wire   [136:0] zext_ln15_1_fu_404_p1;
    reg   [136:0] zext_ln15_1_reg_656;
    wire   [0:0] tmp_22_fu_418_p3;
    reg   [0:0] tmp_22_reg_661;
    wire   [136:0] zext_ln18_1_fu_448_p1;
    reg   [136:0] zext_ln18_1_reg_666;
    reg   [31:0] tmp_14_reg_671;
    reg   [0:0] tmp_23_reg_676;
    reg   [0:0] tmp_23_reg_676_pp0_iter1_reg;
    wire   [31:0] val_1_fu_490_p3;
    reg   [31:0] val_1_reg_680;
    wire    ap_CS_fsm_pp0_stage24;
    wire    ap_block_pp0_stage24_11001;
    wire   [0:0] and_ln61_fu_518_p2;
    reg   [0:0] and_ln61_reg_686;
    wire    ap_CS_fsm_pp0_stage25;
    wire    ap_block_pp0_stage25_11001;
    reg   [0:0] and_ln61_reg_686_pp0_iter1_reg;
    wire   [6:0] trunc_ln62_1_fu_531_p1;
    reg   [6:0] trunc_ln62_1_reg_695;
    wire    ap_block_pp0_stage27_11001;
    reg   [13:0] ogm_grid_addr_reg_705;
    wire    ap_CS_fsm_pp0_stage28;
    wire    ap_block_pp0_stage28_11001;
    reg   [63:0] ogm_grid_load_reg_710;
    wire    ap_CS_fsm_pp0_stage29;
    wire    ap_block_pp0_stage29_11001;
    reg   [63:0] mul17_i_reg_716;
    wire    ap_CS_fsm_pp0_stage36;
    wire    ap_block_pp0_stage36_11001;
    reg   [63:0] sub23_i_reg_721;
    reg   [63:0] div_i_reg_726;
    wire    ap_CS_fsm_pp0_stage26;
    wire    ap_block_pp0_stage26_11001;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire   [63:0] zext_ln62_2_fu_538_p1;
    wire    ap_block_pp0_stage28;
    reg   [31:0] i_fu_82;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    wire    ap_loop_init;
    reg   [31:0] ap_sig_allocacmp_i_4;
    wire    ap_block_pp0_stage0;
    wire    ap_block_pp0_stage27;
    reg   [63:0] grp_fu_129_p0;
    reg   [63:0] grp_fu_129_p1;
    wire    ap_block_pp0_stage14;
    wire    ap_CS_fsm_pp0_stage15;
    wire    ap_block_pp0_stage15;
    wire    ap_CS_fsm_pp0_stage30;
    wire    ap_block_pp0_stage30;
    reg   [63:0] grp_fu_135_p0;
    reg   [63:0] grp_fu_135_p1;
    wire    ap_block_pp0_stage7;
    wire    ap_block_pp0_stage8;
    wire    ap_block_pp0_stage37;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6;
    wire   [63:0] bitcast_ln57_fu_182_p1;
    wire   [10:0] tmp_fu_185_p4;
    wire   [51:0] trunc_ln57_fu_195_p1;
    wire   [0:0] icmp_ln57_1_fu_205_p2;
    wire   [0:0] icmp_ln57_fu_199_p2;
    wire   [0:0] or_ln57_fu_211_p2;
    wire   [0:0] or_ln57_1_fu_217_p2;
    wire   [0:0] and_ln57_fu_221_p2;
    wire   [0:0] grp_fu_144_p2;
    wire    ap_block_pp0_stage21;
    wire   [63:0] data_fu_237_p1;
    wire   [51:0] trunc_ln505_fu_259_p1;
    wire   [53:0] mantissa_fu_263_p4;
    wire   [10:0] xs_exp_fu_249_p4;
    wire   [11:0] zext_ln486_fu_277_p1;
    wire   [11:0] add_ln486_fu_281_p2;
    wire   [10:0] sub_ln18_fu_295_p2;
    wire  signed [11:0] sext_ln18_fu_301_p1;
    wire   [11:0] select_ln18_fu_305_p3;
    wire  signed [31:0] sext_ln18_1_fu_313_p1;
    wire   [136:0] lshr_ln18_fu_321_p2;
    wire    ap_block_pp0_stage22;
    wire   [136:0] shl_ln18_fu_337_p2;
    wire   [31:0] tmp_13_fu_341_p4;
    wire    ap_block_pp0_stage23;
    wire   [31:0] result_1_fu_357_p2;
    wire   [63:0] data_2_fu_368_p1;
    wire   [51:0] trunc_ln505_1_fu_390_p1;
    wire   [53:0] mantissa_1_fu_394_p4;
    wire   [10:0] xs_exp_1_fu_380_p4;
    wire   [11:0] zext_ln486_1_fu_408_p1;
    wire   [11:0] add_ln486_1_fu_412_p2;
    wire   [10:0] sub_ln18_1_fu_426_p2;
    wire  signed [11:0] sext_ln18_2_fu_432_p1;
    wire   [11:0] select_ln18_2_fu_436_p3;
    wire  signed [31:0] sext_ln18_3_fu_444_p1;
    wire   [136:0] lshr_ln18_1_fu_452_p2;
    wire    ap_block_pp0_stage24;
    wire   [136:0] shl_ln18_1_fu_476_p2;
    wire   [31:0] tmp_15_fu_480_p4;
    wire    ap_block_pp0_stage25;
    wire   [31:0] result_4_fu_496_p2;
    wire   [31:0] result_6_fu_501_p3;
    wire   [0:0] icmp_ln61_1_fu_512_p2;
    wire   [0:0] icmp_ln61_fu_507_p2;
    wire   [6:0] trunc_ln62_fu_524_p1;
    wire   [13:0] grp_fu_542_p3;
    wire   [6:0] grp_fu_542_p0;
    wire   [6:0] grp_fu_542_p1;
    wire   [6:0] grp_fu_542_p2;
    reg   [1:0] grp_fu_129_opcode;
    wire    ap_block_pp0_stage14_00001;
    wire    ap_block_pp0_stage15_00001;
    wire    ap_block_pp0_stage30_00001;
    wire    ap_block_pp0_stage6_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [68:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to1;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_block_pp0_stage13_subdone;
    wire    ap_block_pp0_stage14_subdone;
    wire    ap_block_pp0_stage15_subdone;
    wire    ap_block_pp0_stage16_subdone;
    wire    ap_block_pp0_stage17_subdone;
    wire    ap_block_pp0_stage18_subdone;
    wire    ap_block_pp0_stage19_subdone;
    wire    ap_block_pp0_stage20_subdone;
    wire    ap_block_pp0_stage21_subdone;
    wire    ap_block_pp0_stage22_subdone;
    wire    ap_block_pp0_stage23_subdone;
    wire    ap_block_pp0_stage24_subdone;
    wire    ap_block_pp0_stage25_subdone;
    wire    ap_block_pp0_stage26_subdone;
    wire    ap_block_pp0_stage28_subdone;
    wire    ap_block_pp0_stage29_subdone;
    wire    ap_block_pp0_stage30_subdone;
    wire    ap_block_pp0_stage31_subdone;
    wire    ap_block_pp0_stage32_subdone;
    wire    ap_block_pp0_stage33_subdone;
    wire    ap_block_pp0_stage34_subdone;
    wire    ap_block_pp0_stage35_subdone;
    wire    ap_block_pp0_stage36_subdone;
    wire    ap_block_pp0_stage37_subdone;
    wire    ap_block_pp0_stage38_subdone;
    wire    ap_block_pp0_stage39_subdone;
    wire    ap_block_pp0_stage40_subdone;
    wire    ap_block_pp0_stage41_subdone;
    wire    ap_block_pp0_stage42_subdone;
    wire    ap_block_pp0_stage43_subdone;
    wire    ap_block_pp0_stage44_subdone;
    wire    ap_block_pp0_stage45_subdone;
    wire    ap_block_pp0_stage46_subdone;
    wire    ap_block_pp0_stage47_subdone;
    wire    ap_block_pp0_stage48_subdone;
    wire    ap_block_pp0_stage49_subdone;
    wire    ap_block_pp0_stage50_subdone;
    wire    ap_block_pp0_stage51_subdone;
    wire    ap_block_pp0_stage52_subdone;
    wire    ap_block_pp0_stage53_subdone;
    wire    ap_block_pp0_stage54_subdone;
    wire    ap_block_pp0_stage55_subdone;
    wire    ap_block_pp0_stage56_subdone;
    wire    ap_block_pp0_stage57_subdone;
    wire    ap_block_pp0_stage58_subdone;
    wire    ap_block_pp0_stage59_subdone;
    wire    ap_block_pp0_stage60_subdone;
    wire    ap_block_pp0_stage61_subdone;
    wire    ap_block_pp0_stage62_subdone;
    wire    ap_block_pp0_stage63_subdone;
    wire    ap_block_pp0_stage64_subdone;
    wire    ap_block_pp0_stage65_subdone;
    wire    ap_block_pp0_stage66_subdone;
    wire    ap_block_pp0_stage67_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire   [13:0] grp_fu_542_p00;
    wire   [13:0] grp_fu_542_p20;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 69'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 i_fu_82 = 32'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U66 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_135_p0),
        .din1(grp_fu_135_p1),
        .ce(1'b1),
        .dout(grp_fu_135_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_U68 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(conv_i_reg_593),
        .din1(measurement),
        .ce(1'b1),
        .opcode(5'd4),
        .dout(grp_fu_144_p2)
    );

    main_sitodp_32ns_64_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) sitodp_32ns_64_6_no_dsp_1_U69 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(ap_sig_allocacmp_i_4),
        .ce(1'b1),
        .dout(grp_fu_148_p1)
    );

    main_mac_muladd_7ns_7ns_7ns_14_4_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(7),
        .din1_WIDTH(7),
        .din2_WIDTH(7),
        .dout_WIDTH(14)
    ) mac_muladd_7ns_7ns_7ns_14_4_1_U70 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_542_p0),
        .din1(grp_fu_542_p1),
        .din2(grp_fu_542_p2),
        .ce(1'b1),
        .dout(grp_fu_542_p3)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage27),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage27) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage27_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage27)) begin
                ap_enable_reg_pp0_iter0_reg <= 1'b0;
            end else if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (1'b0 == ap_block_pp0_stage27_subdone))) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage68) & (1'b0 == ap_block_pp0_stage68_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            i_fu_82 <= 32'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'd1 == and_ln57_1_reg_600) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8_11001))) begin
            i_fu_82 <= i_5_reg_588;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7_11001))) begin
            and_ln57_1_reg_600 <= and_ln57_1_fu_227_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage25) & (1'b0 == ap_block_pp0_stage25_11001))) begin
            and_ln61_reg_686 <= and_ln61_fu_518_p2;
            and_ln61_reg_686_pp0_iter1_reg <= and_ln61_reg_686;
            trunc_ln62_1_reg_695 <= trunc_ln62_1_fu_531_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5_11001))) begin
            conv_i_reg_593 <= grp_fu_148_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage26) & (1'b0 == ap_block_pp0_stage26_11001))) begin
            div_i_reg_726 <= grp_fu_194_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            i_5_reg_588 <= i_5_fu_176_p2;
            icmp_ln57_2_reg_578 <= icmp_ln57_2_fu_164_p2;
            icmp_ln57_3_reg_583 <= icmp_ln57_3_fu_170_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36) & (1'b0 == ap_block_pp0_stage36_11001))) begin
            mul17_i_reg_716 <= grp_fu_135_p2;
            sub23_i_reg_721 <= grp_fu_172_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_11001))) begin
            mul5_i_reg_609 <= grp_fu_135_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13) & (1'b0 == ap_block_pp0_stage13_11001))) begin
            mul_i_reg_604 <= grp_fu_135_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28_11001))) begin
            ogm_grid_addr_reg_705 <= zext_ln62_2_fu_538_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29) & (1'b0 == ap_block_pp0_stage29_11001))) begin
            ogm_grid_load_reg_710 <= ogm_grid_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20) & (1'b0 == ap_block_pp0_stage20_11001)))) begin
            reg_151 <= grp_fu_172_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage23) & (1'b0 == ap_block_pp0_stage23_11001))) begin
            result_reg_645 <= result_fu_362_p3;
            tmp_14_reg_671 <= {{lshr_ln18_1_fu_452_p2[84:53]}};
            tmp_22_reg_661 <= add_ln486_1_fu_412_p2[32'd11];
            tmp_23_reg_676 <= result_fu_362_p3[32'd31];
            tmp_23_reg_676_pp0_iter1_reg <= tmp_23_reg_676;
            xs_sign_1_reg_651 <= data_2_fu_368_p1[32'd63];
            zext_ln15_1_reg_656[52 : 1] <= zext_ln15_1_fu_404_p1[52 : 1];
            zext_ln18_1_reg_666[31 : 0] <= zext_ln18_1_fu_448_p1[31 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage21) & (1'b0 == ap_block_pp0_stage21_11001))) begin
            tmp_20_reg_624 <= add_ln486_fu_281_p2[32'd11];
            tmp_s_reg_634 <= {{lshr_ln18_fu_321_p2[84:53]}};
            xs_sign_reg_614 <= data_fu_237_p1[32'd63];
            zext_ln15_reg_619[52 : 1] <= zext_ln15_fu_273_p1[52 : 1];
            zext_ln18_reg_629[31 : 0] <= zext_ln18_fu_317_p1[31 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage24) & (1'b0 == ap_block_pp0_stage24_11001))) begin
            val_1_reg_680 <= val_1_fu_490_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage22) & (1'b0 == ap_block_pp0_stage22_11001))) begin
            val_reg_639 <= val_fu_351_p3;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (1'd0 == and_ln57_1_reg_600) & (1'b0 == ap_block_pp0_stage27_subdone))) begin
            ap_condition_exit_pp0_iter0_stage27 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage27 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage27) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage27_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b0)) begin
            ap_idle_pp0_1to1 = 1'b1;
        end else begin
            ap_idle_pp0_1to1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage68) & (1'b0 == ap_block_pp0_stage68_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_i_4 = 32'd0;
        end else begin
            ap_sig_allocacmp_i_4 = i_fu_82;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'd1 == and_ln61_reg_686) & (1'd1 == and_ln57_1_reg_600) & (tmp_23_reg_676 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30_00001))) begin
            grp_fu_129_opcode = 2'd1;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'd1 == and_ln57_1_reg_600) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15_00001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'd1 == and_ln57_1_reg_600) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14_00001)))) begin
            grp_fu_129_opcode = 2'd0;
        end else begin
            grp_fu_129_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
                grp_fu_129_p0 = 64'd4607182418800017408;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15))) begin
                grp_fu_129_p0 = mul5_i_reg_609;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14))) begin
                grp_fu_129_p0 = mul_i_reg_604;
            end else begin
                grp_fu_129_p0 = 'bx;
            end
        end else begin
            grp_fu_129_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_129_p1 = ogm_grid_load_reg_710;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15) & (1'b0 == ap_block_pp0_stage15)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14) & (1'b0 == ap_block_pp0_stage14)))) begin
            grp_fu_129_p1 = 64'd4632233691727265792;
        end else begin
            grp_fu_129_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
            grp_fu_135_p0 = ogm_grid_load_reg_710;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7)))) begin
            grp_fu_135_p0 = conv_i_reg_593;
        end else begin
            grp_fu_135_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b1 == ap_CS_fsm_pp0_stage30) & (1'b0 == ap_block_pp0_stage30))) begin
                grp_fu_135_p1 = 64'd4599075939470750516;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage8) & (1'b0 == ap_block_pp0_stage8))) begin
                grp_fu_135_p1 = dy;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage7) & (1'b0 == ap_block_pp0_stage7))) begin
                grp_fu_135_p1 = dx;
            end else begin
                grp_fu_135_p1 = 'bx;
            end
        end else begin
            grp_fu_135_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (1'b0 == ap_block_pp0_stage27))) begin
            ogm_grid_address0 = ogm_grid_addr_reg_705;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28))) begin
            ogm_grid_address0 = zext_ln62_2_fu_538_p1;
        end else begin
            ogm_grid_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27) & (1'b0 == ap_block_pp0_stage27_11001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28) & (1'b0 == ap_block_pp0_stage28_11001)))) begin
            ogm_grid_ce0 = 1'b1;
        end else begin
            ogm_grid_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'd1 == and_ln61_reg_686_pp0_iter1_reg) & (tmp_23_reg_676_pp0_iter1_reg == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage27) & (1'b0 == ap_block_pp0_stage27_11001))) begin
            ogm_grid_we0 = 1'b1;
        end else begin
            ogm_grid_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_idle_pp0_1to1 == 1'b1) & (ap_start_int == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            ap_ST_fsm_pp0_stage14: begin
                if ((1'b0 == ap_block_pp0_stage14_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end
            end
            ap_ST_fsm_pp0_stage15: begin
                if ((1'b0 == ap_block_pp0_stage15_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end
            end
            ap_ST_fsm_pp0_stage16: begin
                if ((1'b0 == ap_block_pp0_stage16_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end
            end
            ap_ST_fsm_pp0_stage17: begin
                if ((1'b0 == ap_block_pp0_stage17_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end
            end
            ap_ST_fsm_pp0_stage18: begin
                if ((1'b0 == ap_block_pp0_stage18_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end
            end
            ap_ST_fsm_pp0_stage19: begin
                if ((1'b0 == ap_block_pp0_stage19_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end
            end
            ap_ST_fsm_pp0_stage20: begin
                if ((1'b0 == ap_block_pp0_stage20_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end
            end
            ap_ST_fsm_pp0_stage21: begin
                if ((1'b0 == ap_block_pp0_stage21_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end
            end
            ap_ST_fsm_pp0_stage22: begin
                if ((1'b0 == ap_block_pp0_stage22_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end
            end
            ap_ST_fsm_pp0_stage23: begin
                if ((1'b0 == ap_block_pp0_stage23_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end
            end
            ap_ST_fsm_pp0_stage24: begin
                if ((1'b0 == ap_block_pp0_stage24_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end
            end
            ap_ST_fsm_pp0_stage25: begin
                if ((1'b0 == ap_block_pp0_stage25_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end
            end
            ap_ST_fsm_pp0_stage26: begin
                if ((1'b0 == ap_block_pp0_stage26_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end
            end
            ap_ST_fsm_pp0_stage27: begin
                if ((1'b1 == ap_condition_exit_pp0_iter0_stage27)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage27_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end
            end
            ap_ST_fsm_pp0_stage28: begin
                if ((1'b0 == ap_block_pp0_stage28_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end
            end
            ap_ST_fsm_pp0_stage29: begin
                if ((1'b0 == ap_block_pp0_stage29_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end
            end
            ap_ST_fsm_pp0_stage30: begin
                if ((1'b0 == ap_block_pp0_stage30_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end
            end
            ap_ST_fsm_pp0_stage31: begin
                if ((1'b0 == ap_block_pp0_stage31_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end
            end
            ap_ST_fsm_pp0_stage32: begin
                if ((1'b0 == ap_block_pp0_stage32_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end
            end
            ap_ST_fsm_pp0_stage33: begin
                if ((1'b0 == ap_block_pp0_stage33_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end
            end
            ap_ST_fsm_pp0_stage34: begin
                if ((1'b0 == ap_block_pp0_stage34_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end
            end
            ap_ST_fsm_pp0_stage35: begin
                if ((1'b0 == ap_block_pp0_stage35_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end
            end
            ap_ST_fsm_pp0_stage36: begin
                if ((1'b0 == ap_block_pp0_stage36_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end
            end
            ap_ST_fsm_pp0_stage37: begin
                if ((1'b0 == ap_block_pp0_stage37_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end
            end
            ap_ST_fsm_pp0_stage38: begin
                if ((1'b0 == ap_block_pp0_stage38_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end
            end
            ap_ST_fsm_pp0_stage39: begin
                if ((1'b0 == ap_block_pp0_stage39_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end
            end
            ap_ST_fsm_pp0_stage40: begin
                if ((1'b0 == ap_block_pp0_stage40_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end
            end
            ap_ST_fsm_pp0_stage41: begin
                if ((1'b0 == ap_block_pp0_stage41_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end
            end
            ap_ST_fsm_pp0_stage42: begin
                if ((1'b0 == ap_block_pp0_stage42_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end
            end
            ap_ST_fsm_pp0_stage43: begin
                if ((1'b0 == ap_block_pp0_stage43_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end
            end
            ap_ST_fsm_pp0_stage44: begin
                if ((1'b0 == ap_block_pp0_stage44_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end
            end
            ap_ST_fsm_pp0_stage45: begin
                if ((1'b0 == ap_block_pp0_stage45_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end
            end
            ap_ST_fsm_pp0_stage46: begin
                if ((1'b0 == ap_block_pp0_stage46_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end
            end
            ap_ST_fsm_pp0_stage47: begin
                if ((1'b0 == ap_block_pp0_stage47_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end
            end
            ap_ST_fsm_pp0_stage48: begin
                if ((1'b0 == ap_block_pp0_stage48_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end
            end
            ap_ST_fsm_pp0_stage49: begin
                if ((1'b0 == ap_block_pp0_stage49_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end
            end
            ap_ST_fsm_pp0_stage50: begin
                if ((1'b0 == ap_block_pp0_stage50_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end
            end
            ap_ST_fsm_pp0_stage51: begin
                if ((1'b0 == ap_block_pp0_stage51_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end
            end
            ap_ST_fsm_pp0_stage52: begin
                if ((1'b0 == ap_block_pp0_stage52_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end
            end
            ap_ST_fsm_pp0_stage53: begin
                if ((1'b0 == ap_block_pp0_stage53_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end
            end
            ap_ST_fsm_pp0_stage54: begin
                if ((1'b0 == ap_block_pp0_stage54_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end
            end
            ap_ST_fsm_pp0_stage55: begin
                if ((1'b0 == ap_block_pp0_stage55_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end
            end
            ap_ST_fsm_pp0_stage56: begin
                if ((1'b0 == ap_block_pp0_stage56_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end
            end
            ap_ST_fsm_pp0_stage57: begin
                if ((1'b0 == ap_block_pp0_stage57_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end
            end
            ap_ST_fsm_pp0_stage58: begin
                if ((1'b0 == ap_block_pp0_stage58_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end
            end
            ap_ST_fsm_pp0_stage59: begin
                if ((1'b0 == ap_block_pp0_stage59_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end
            end
            ap_ST_fsm_pp0_stage60: begin
                if ((1'b0 == ap_block_pp0_stage60_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end
            end
            ap_ST_fsm_pp0_stage61: begin
                if ((1'b0 == ap_block_pp0_stage61_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end
            end
            ap_ST_fsm_pp0_stage62: begin
                if ((1'b0 == ap_block_pp0_stage62_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end
            end
            ap_ST_fsm_pp0_stage63: begin
                if ((1'b0 == ap_block_pp0_stage63_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end
            end
            ap_ST_fsm_pp0_stage64: begin
                if ((1'b0 == ap_block_pp0_stage64_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end
            end
            ap_ST_fsm_pp0_stage65: begin
                if ((1'b0 == ap_block_pp0_stage65_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end
            end
            ap_ST_fsm_pp0_stage66: begin
                if ((1'b0 == ap_block_pp0_stage66_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end
            end
            ap_ST_fsm_pp0_stage67: begin
                if ((1'b0 == ap_block_pp0_stage67_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end
            end
            ap_ST_fsm_pp0_stage68: begin
                if ((1'b0 == ap_block_pp0_stage68_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln486_1_fu_412_p2 = ($signed(zext_ln486_1_fu_408_p1) + $signed(12'd3073));

    assign add_ln486_fu_281_p2 = ($signed(zext_ln486_fu_277_p1) + $signed(12'd3073));

    assign and_ln57_1_fu_227_p2 = (grp_fu_144_p2 & and_ln57_fu_221_p2);

    assign and_ln57_fu_221_p2 = (or_ln57_fu_211_p2 & or_ln57_1_fu_217_p2);

    assign and_ln61_fu_518_p2 = (icmp_ln61_fu_507_p2 & icmp_ln61_1_fu_512_p2);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage14 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_pp0_stage15 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_pp0_stage20 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_pp0_stage21 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_pp0_stage22 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_pp0_stage23 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_pp0_stage24 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_pp0_stage25 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_pp0_stage26 = ap_CS_fsm[32'd26];

    assign ap_CS_fsm_pp0_stage27 = ap_CS_fsm[32'd27];

    assign ap_CS_fsm_pp0_stage28 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_pp0_stage29 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_pp0_stage30 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_pp0_stage36 = ap_CS_fsm[32'd36];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage68 = ap_CS_fsm[32'd68];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage53_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage54_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage55_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage56_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage57_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage58_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage59_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage60_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage61_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage62_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage63_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage64_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage65_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage66_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage67_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage68_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage27;

    assign bitcast_ln57_fu_182_p1 = conv_i_reg_593;

    assign data_2_fu_368_p1 = reg_151;

    assign data_fu_237_p1 = reg_151;

    assign grp_fu_172_p_ce = 1'b1;

    assign grp_fu_172_p_din0 = grp_fu_129_p0;

    assign grp_fu_172_p_din1 = grp_fu_129_p1;

    assign grp_fu_172_p_opcode = grp_fu_129_opcode;

    assign grp_fu_194_p_ce = 1'b1;

    assign grp_fu_194_p_din0 = mul17_i_reg_716;

    assign grp_fu_194_p_din1 = sub23_i_reg_721;

    assign grp_fu_542_p0 = grp_fu_542_p00;

    assign grp_fu_542_p00 = trunc_ln62_fu_524_p1;

    assign grp_fu_542_p1 = 14'd100;

    assign grp_fu_542_p2 = grp_fu_542_p20;

    assign grp_fu_542_p20 = trunc_ln62_1_reg_695;

    assign i_5_fu_176_p2 = (ap_sig_allocacmp_i_4 + 32'd1);

    assign icmp_ln57_1_fu_205_p2 = ((trunc_ln57_fu_195_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln57_2_fu_164_p2 = ((tmp_3 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln57_3_fu_170_p2 = ((empty == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln57_fu_199_p2 = ((tmp_fu_185_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln61_1_fu_512_p2 = ((result_6_fu_501_p3 < 32'd100) ? 1'b1 : 1'b0);

    assign icmp_ln61_fu_507_p2 = (($signed(result_reg_645) < $signed(32'd100)) ? 1'b1 : 1'b0);

    assign lshr_ln18_1_fu_452_p2 = zext_ln15_1_fu_404_p1 >> zext_ln18_1_fu_448_p1;

    assign lshr_ln18_fu_321_p2 = zext_ln15_fu_273_p1 >> zext_ln18_fu_317_p1;

    assign mantissa_1_fu_394_p4 = {{{{1'd1}, {trunc_ln505_1_fu_390_p1}}}, {1'd0}};

    assign mantissa_fu_263_p4 = {{{{1'd1}, {trunc_ln505_fu_259_p1}}}, {1'd0}};

    assign ogm_grid_d0 = div_i_reg_726;

    assign or_ln57_1_fu_217_p2 = (icmp_ln57_3_reg_583 | icmp_ln57_2_reg_578);

    assign or_ln57_fu_211_p2 = (icmp_ln57_fu_199_p2 | icmp_ln57_1_fu_205_p2);

    assign result_1_fu_357_p2 = (32'd0 - val_reg_639);

    assign result_4_fu_496_p2 = (32'd0 - val_1_reg_680);

    assign result_6_fu_501_p3 = ((xs_sign_1_reg_651[0:0] == 1'b1) ? result_4_fu_496_p2 : val_1_reg_680);

    assign result_fu_362_p3 = ((xs_sign_reg_614[0:0] == 1'b1) ? result_1_fu_357_p2 : val_reg_639);

    assign select_ln18_2_fu_436_p3 = ((tmp_22_fu_418_p3[0:0] == 1'b1) ? sext_ln18_2_fu_432_p1 : add_ln486_1_fu_412_p2);

    assign select_ln18_fu_305_p3 = ((tmp_20_fu_287_p3[0:0] == 1'b1) ? sext_ln18_fu_301_p1 : add_ln486_fu_281_p2);

    assign sext_ln18_1_fu_313_p1 = $signed(select_ln18_fu_305_p3);

    assign sext_ln18_2_fu_432_p1 = $signed(sub_ln18_1_fu_426_p2);

    assign sext_ln18_3_fu_444_p1 = $signed(select_ln18_2_fu_436_p3);

    assign sext_ln18_fu_301_p1 = $signed(sub_ln18_fu_295_p2);

    assign shl_ln18_1_fu_476_p2 = zext_ln15_1_reg_656 << zext_ln18_1_reg_666;

    assign shl_ln18_fu_337_p2 = zext_ln15_reg_619 << zext_ln18_reg_629;

    assign sub_ln18_1_fu_426_p2 = (11'd1023 - xs_exp_1_fu_380_p4);

    assign sub_ln18_fu_295_p2 = (11'd1023 - xs_exp_fu_249_p4);

    assign tmp_13_fu_341_p4 = {{shl_ln18_fu_337_p2[84:53]}};

    assign tmp_15_fu_480_p4 = {{shl_ln18_1_fu_476_p2[84:53]}};

    assign tmp_20_fu_287_p3 = add_ln486_fu_281_p2[32'd11];

    assign tmp_22_fu_418_p3 = add_ln486_1_fu_412_p2[32'd11];

    assign tmp_fu_185_p4 = {{bitcast_ln57_fu_182_p1[62:52]}};

    assign trunc_ln505_1_fu_390_p1 = data_2_fu_368_p1[51:0];

    assign trunc_ln505_fu_259_p1 = data_fu_237_p1[51:0];

    assign trunc_ln57_fu_195_p1 = bitcast_ln57_fu_182_p1[51:0];

    assign trunc_ln62_1_fu_531_p1 = result_6_fu_501_p3[6:0];

    assign trunc_ln62_fu_524_p1 = result_reg_645[6:0];

    assign val_1_fu_490_p3 = ((tmp_22_reg_661[0:0] == 1'b1) ? tmp_14_reg_671 : tmp_15_fu_480_p4);

    assign val_fu_351_p3 = ((tmp_20_reg_624[0:0] == 1'b1) ? tmp_s_reg_634 : tmp_13_fu_341_p4);

    assign xs_exp_1_fu_380_p4 = {{data_2_fu_368_p1[62:52]}};

    assign xs_exp_fu_249_p4 = {{data_fu_237_p1[62:52]}};

    assign zext_ln15_1_fu_404_p1 = mantissa_1_fu_394_p4;

    assign zext_ln15_fu_273_p1 = mantissa_fu_263_p4;

    assign zext_ln18_1_fu_448_p1 = $unsigned(sext_ln18_3_fu_444_p1);

    assign zext_ln18_fu_317_p1 = $unsigned(sext_ln18_1_fu_313_p1);

    assign zext_ln486_1_fu_408_p1 = xs_exp_1_fu_380_p4;

    assign zext_ln486_fu_277_p1 = xs_exp_fu_249_p4;

    assign zext_ln62_2_fu_538_p1 = grp_fu_542_p3;

    always @(posedge ap_clk) begin
        zext_ln15_reg_619[0] <= 1'b0;
        zext_ln15_reg_619[136:53] <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        zext_ln18_reg_629[136:32] <= 105'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        zext_ln15_1_reg_656[0] <= 1'b0;
        zext_ln15_1_reg_656[136:53] <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        zext_ln18_1_reg_666[136:32] <= 105'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_main_Pipeline_VITIS_LOOP_57_1
