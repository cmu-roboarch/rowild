/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_3 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    empty,
    l_cAxes_address0,
    l_cAxes_ce0,
    l_cAxes_we0,
    l_cAxes_d0
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [4:0] empty;
    output [5:0] l_cAxes_address0;
    output l_cAxes_ce0;
    output l_cAxes_we0;
    output [63:0] l_cAxes_d0;

    reg ap_idle;
    reg l_cAxes_ce0;
    reg l_cAxes_we0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] exitcond227_fu_98_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire   [5:0] empty_68_fu_133_p2;
    reg   [5:0] empty_68_reg_226;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] p_cast1_fu_192_p1;
    wire    ap_block_pp0_stage0;
    reg   [3:0] phi_urem9_fu_44;
    wire   [3:0] idx_urem11_fu_164_p3;
    wire    ap_loop_init;
    reg   [7:0] phi_mul7_fu_48;
    wire   [7:0] next_mul8_fu_113_p2;
    reg   [7:0] ap_sig_allocacmp_phi_mul7_load;
    reg   [3:0] empty_65_fu_52;
    wire   [3:0] empty_66_fu_104_p2;
    reg   [3:0] ap_sig_allocacmp_p_load;
    wire   [1:0] tmp_21_fu_119_p4;
    wire  signed [5:0] p_cast_fu_76_p1;
    wire   [5:0] tmp_42_cast_fu_129_p1;
    wire   [3:0] next_urem10_fu_152_p2;
    wire   [0:0] empty_67_fu_158_p2;
    wire   [5:0] empty_69_fu_172_p2;
    wire   [5:0] empty_70_fu_177_p2;
    wire   [5:0] phi_urem9_cast_fu_182_p1;
    wire   [5:0] empty_71_fu_186_p2;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 phi_urem9_fu_44 = 4'd0;
        #0 phi_mul7_fu_48 = 8'd0;
        #0 empty_65_fu_52 = 4'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((exitcond227_fu_98_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                empty_65_fu_52 <= empty_66_fu_104_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                empty_65_fu_52 <= 4'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((exitcond227_fu_98_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                phi_mul7_fu_48 <= next_mul8_fu_113_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                phi_mul7_fu_48 <= 8'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                phi_urem9_fu_44 <= 4'd0;
            end else if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
                phi_urem9_fu_44 <= idx_urem11_fu_164_p3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            empty_68_reg_226 <= empty_68_fu_133_p2;
        end
    end

    always @(*) begin
        if (((exitcond227_fu_98_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_p_load = 4'd0;
        end else begin
            ap_sig_allocacmp_p_load = empty_65_fu_52;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_phi_mul7_load = 8'd0;
        end else begin
            ap_sig_allocacmp_phi_mul7_load = phi_mul7_fu_48;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_cAxes_ce0 = 1'b1;
        end else begin
            l_cAxes_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_cAxes_we0 = 1'b1;
        end else begin
            l_cAxes_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign empty_66_fu_104_p2 = (ap_sig_allocacmp_p_load + 4'd1);

    assign empty_67_fu_158_p2 = ((next_urem10_fu_152_p2 < 4'd3) ? 1'b1 : 1'b0);

    assign empty_68_fu_133_p2 = ($signed(p_cast_fu_76_p1) + $signed(tmp_42_cast_fu_129_p1));

    assign empty_69_fu_172_p2 = empty_68_reg_226 << 6'd2;

    assign empty_70_fu_177_p2 = (empty_69_fu_172_p2 - empty_68_reg_226);

    assign empty_71_fu_186_p2 = (empty_70_fu_177_p2 + phi_urem9_cast_fu_182_p1);

    assign exitcond227_fu_98_p2 = ((ap_sig_allocacmp_p_load == 4'd9) ? 1'b1 : 1'b0);

    assign idx_urem11_fu_164_p3 = ((empty_67_fu_158_p2[0:0] == 1'b1) ? next_urem10_fu_152_p2 : 4'd0);

    assign l_cAxes_address0 = p_cast1_fu_192_p1;

    assign l_cAxes_d0 = 64'd0;

    assign next_mul8_fu_113_p2 = (ap_sig_allocacmp_phi_mul7_load + 8'd22);

    assign next_urem10_fu_152_p2 = (phi_urem9_fu_44 + 4'd1);

    assign p_cast1_fu_192_p1 = empty_71_fu_186_p2;

    assign p_cast_fu_76_p1 = $signed(empty);

    assign phi_urem9_cast_fu_182_p1 = phi_urem9_fu_44;

    assign tmp_21_fu_119_p4 = {{ap_sig_allocacmp_phi_mul7_load[7:6]}};

    assign tmp_42_cast_fu_129_p1 = tmp_21_fu_119_p4;

endmodule  //main_main_Pipeline_3
