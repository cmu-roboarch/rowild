/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_cuboidCuboidCollision_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    axes1_address0,
    axes1_ce0,
    axes1_q0,
    axes1_address1,
    axes1_ce1,
    axes1_q1,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    axes2_address0,
    axes2_ce0,
    axes2_q0,
    axes2_address1,
    axes2_ce1,
    axes2_q1,
    ap_return,
    grp_fu_1754_p_din0,
    grp_fu_1754_p_din1,
    grp_fu_1754_p_opcode,
    grp_fu_1754_p_dout0,
    grp_fu_1754_p_ce,
    grp_fu_1762_p_din0,
    grp_fu_1762_p_din1,
    grp_fu_1762_p_opcode,
    grp_fu_1762_p_dout0,
    grp_fu_1762_p_ce,
    grp_fu_1766_p_din0,
    grp_fu_1766_p_din1,
    grp_fu_1766_p_opcode,
    grp_fu_1766_p_dout0,
    grp_fu_1766_p_ce,
    grp_fu_1770_p_din0,
    grp_fu_1770_p_din1,
    grp_fu_1770_p_opcode,
    grp_fu_1770_p_dout0,
    grp_fu_1770_p_ce,
    grp_fu_1774_p_din0,
    grp_fu_1774_p_din1,
    grp_fu_1774_p_opcode,
    grp_fu_1774_p_dout0,
    grp_fu_1774_p_ce,
    grp_fu_1778_p_din0,
    grp_fu_1778_p_din1,
    grp_fu_1778_p_opcode,
    grp_fu_1778_p_dout0,
    grp_fu_1778_p_ce,
    grp_fu_1758_p_din0,
    grp_fu_1758_p_din1,
    grp_fu_1758_p_dout0,
    grp_fu_1758_p_ce,
    grp_fu_1782_p_din0,
    grp_fu_1782_p_din1,
    grp_fu_1782_p_dout0,
    grp_fu_1782_p_ce,
    grp_fu_1786_p_din0,
    grp_fu_1786_p_din1,
    grp_fu_1786_p_dout0,
    grp_fu_1786_p_ce,
    grp_fu_1790_p_din0,
    grp_fu_1790_p_din1,
    grp_fu_1790_p_dout0,
    grp_fu_1790_p_ce,
    grp_fu_1794_p_din0,
    grp_fu_1794_p_din1,
    grp_fu_1794_p_opcode,
    grp_fu_1794_p_dout0,
    grp_fu_1794_p_ce,
    grp_fu_1798_p_din0,
    grp_fu_1798_p_din1,
    grp_fu_1798_p_dout0,
    grp_fu_1798_p_ce
);

    parameter ap_ST_fsm_state1 = 104'd1;
    parameter ap_ST_fsm_state2 = 104'd2;
    parameter ap_ST_fsm_state3 = 104'd4;
    parameter ap_ST_fsm_state4 = 104'd8;
    parameter ap_ST_fsm_state5 = 104'd16;
    parameter ap_ST_fsm_state6 = 104'd32;
    parameter ap_ST_fsm_state7 = 104'd64;
    parameter ap_ST_fsm_state8 = 104'd128;
    parameter ap_ST_fsm_state9 = 104'd256;
    parameter ap_ST_fsm_state10 = 104'd512;
    parameter ap_ST_fsm_state11 = 104'd1024;
    parameter ap_ST_fsm_state12 = 104'd2048;
    parameter ap_ST_fsm_state13 = 104'd4096;
    parameter ap_ST_fsm_state14 = 104'd8192;
    parameter ap_ST_fsm_state15 = 104'd16384;
    parameter ap_ST_fsm_state16 = 104'd32768;
    parameter ap_ST_fsm_state17 = 104'd65536;
    parameter ap_ST_fsm_state18 = 104'd131072;
    parameter ap_ST_fsm_state19 = 104'd262144;
    parameter ap_ST_fsm_state20 = 104'd524288;
    parameter ap_ST_fsm_state21 = 104'd1048576;
    parameter ap_ST_fsm_state22 = 104'd2097152;
    parameter ap_ST_fsm_state23 = 104'd4194304;
    parameter ap_ST_fsm_state24 = 104'd8388608;
    parameter ap_ST_fsm_state25 = 104'd16777216;
    parameter ap_ST_fsm_state26 = 104'd33554432;
    parameter ap_ST_fsm_state27 = 104'd67108864;
    parameter ap_ST_fsm_state28 = 104'd134217728;
    parameter ap_ST_fsm_state29 = 104'd268435456;
    parameter ap_ST_fsm_state30 = 104'd536870912;
    parameter ap_ST_fsm_state31 = 104'd1073741824;
    parameter ap_ST_fsm_state32 = 104'd2147483648;
    parameter ap_ST_fsm_state33 = 104'd4294967296;
    parameter ap_ST_fsm_state34 = 104'd8589934592;
    parameter ap_ST_fsm_state35 = 104'd17179869184;
    parameter ap_ST_fsm_state36 = 104'd34359738368;
    parameter ap_ST_fsm_state37 = 104'd68719476736;
    parameter ap_ST_fsm_state38 = 104'd137438953472;
    parameter ap_ST_fsm_state39 = 104'd274877906944;
    parameter ap_ST_fsm_state40 = 104'd549755813888;
    parameter ap_ST_fsm_state41 = 104'd1099511627776;
    parameter ap_ST_fsm_state42 = 104'd2199023255552;
    parameter ap_ST_fsm_state43 = 104'd4398046511104;
    parameter ap_ST_fsm_state44 = 104'd8796093022208;
    parameter ap_ST_fsm_state45 = 104'd17592186044416;
    parameter ap_ST_fsm_state46 = 104'd35184372088832;
    parameter ap_ST_fsm_state47 = 104'd70368744177664;
    parameter ap_ST_fsm_state48 = 104'd140737488355328;
    parameter ap_ST_fsm_state49 = 104'd281474976710656;
    parameter ap_ST_fsm_state50 = 104'd562949953421312;
    parameter ap_ST_fsm_state51 = 104'd1125899906842624;
    parameter ap_ST_fsm_state52 = 104'd2251799813685248;
    parameter ap_ST_fsm_state53 = 104'd4503599627370496;
    parameter ap_ST_fsm_state54 = 104'd9007199254740992;
    parameter ap_ST_fsm_state55 = 104'd18014398509481984;
    parameter ap_ST_fsm_state56 = 104'd36028797018963968;
    parameter ap_ST_fsm_state57 = 104'd72057594037927936;
    parameter ap_ST_fsm_state58 = 104'd144115188075855872;
    parameter ap_ST_fsm_state59 = 104'd288230376151711744;
    parameter ap_ST_fsm_state60 = 104'd576460752303423488;
    parameter ap_ST_fsm_state61 = 104'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 104'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 104'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 104'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 104'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 104'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 104'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 104'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 104'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 104'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 104'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 104'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 104'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 104'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 104'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 104'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 104'd75557863725914323419136;
    parameter ap_ST_fsm_state78 = 104'd151115727451828646838272;
    parameter ap_ST_fsm_state79 = 104'd302231454903657293676544;
    parameter ap_ST_fsm_state80 = 104'd604462909807314587353088;
    parameter ap_ST_fsm_state81 = 104'd1208925819614629174706176;
    parameter ap_ST_fsm_state82 = 104'd2417851639229258349412352;
    parameter ap_ST_fsm_state83 = 104'd4835703278458516698824704;
    parameter ap_ST_fsm_state84 = 104'd9671406556917033397649408;
    parameter ap_ST_fsm_state85 = 104'd19342813113834066795298816;
    parameter ap_ST_fsm_state86 = 104'd38685626227668133590597632;
    parameter ap_ST_fsm_state87 = 104'd77371252455336267181195264;
    parameter ap_ST_fsm_state88 = 104'd154742504910672534362390528;
    parameter ap_ST_fsm_state89 = 104'd309485009821345068724781056;
    parameter ap_ST_fsm_state90 = 104'd618970019642690137449562112;
    parameter ap_ST_fsm_state91 = 104'd1237940039285380274899124224;
    parameter ap_ST_fsm_state92 = 104'd2475880078570760549798248448;
    parameter ap_ST_fsm_state93 = 104'd4951760157141521099596496896;
    parameter ap_ST_fsm_state94 = 104'd9903520314283042199192993792;
    parameter ap_ST_fsm_state95 = 104'd19807040628566084398385987584;
    parameter ap_ST_fsm_state96 = 104'd39614081257132168796771975168;
    parameter ap_ST_fsm_state97 = 104'd79228162514264337593543950336;
    parameter ap_ST_fsm_state98 = 104'd158456325028528675187087900672;
    parameter ap_ST_fsm_state99 = 104'd316912650057057350374175801344;
    parameter ap_ST_fsm_state100 = 104'd633825300114114700748351602688;
    parameter ap_ST_fsm_state101 = 104'd1267650600228229401496703205376;
    parameter ap_ST_fsm_state102 = 104'd2535301200456458802993406410752;
    parameter ap_ST_fsm_state103 = 104'd5070602400912917605986812821504;
    parameter ap_ST_fsm_state104 = 104'd10141204801825835211973625643008;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [5:0] axes1_address0;
    output axes1_ce0;
    input [63:0] axes1_q0;
    output [5:0] axes1_address1;
    output axes1_ce1;
    input [63:0] axes1_q1;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    output [6:0] axes2_address0;
    output axes2_ce0;
    input [63:0] axes2_q0;
    output [6:0] axes2_address1;
    output axes2_ce1;
    input [63:0] axes2_q1;
    output [0:0] ap_return;
    output [63:0] grp_fu_1754_p_din0;
    output [63:0] grp_fu_1754_p_din1;
    output [1:0] grp_fu_1754_p_opcode;
    input [63:0] grp_fu_1754_p_dout0;
    output grp_fu_1754_p_ce;
    output [63:0] grp_fu_1762_p_din0;
    output [63:0] grp_fu_1762_p_din1;
    output [1:0] grp_fu_1762_p_opcode;
    input [63:0] grp_fu_1762_p_dout0;
    output grp_fu_1762_p_ce;
    output [63:0] grp_fu_1766_p_din0;
    output [63:0] grp_fu_1766_p_din1;
    output [1:0] grp_fu_1766_p_opcode;
    input [63:0] grp_fu_1766_p_dout0;
    output grp_fu_1766_p_ce;
    output [63:0] grp_fu_1770_p_din0;
    output [63:0] grp_fu_1770_p_din1;
    output [1:0] grp_fu_1770_p_opcode;
    input [63:0] grp_fu_1770_p_dout0;
    output grp_fu_1770_p_ce;
    output [63:0] grp_fu_1774_p_din0;
    output [63:0] grp_fu_1774_p_din1;
    output [1:0] grp_fu_1774_p_opcode;
    input [63:0] grp_fu_1774_p_dout0;
    output grp_fu_1774_p_ce;
    output [63:0] grp_fu_1778_p_din0;
    output [63:0] grp_fu_1778_p_din1;
    output [1:0] grp_fu_1778_p_opcode;
    input [63:0] grp_fu_1778_p_dout0;
    output grp_fu_1778_p_ce;
    output [63:0] grp_fu_1758_p_din0;
    output [63:0] grp_fu_1758_p_din1;
    input [63:0] grp_fu_1758_p_dout0;
    output grp_fu_1758_p_ce;
    output [63:0] grp_fu_1782_p_din0;
    output [63:0] grp_fu_1782_p_din1;
    input [63:0] grp_fu_1782_p_dout0;
    output grp_fu_1782_p_ce;
    output [63:0] grp_fu_1786_p_din0;
    output [63:0] grp_fu_1786_p_din1;
    input [63:0] grp_fu_1786_p_dout0;
    output grp_fu_1786_p_ce;
    output [63:0] grp_fu_1790_p_din0;
    output [63:0] grp_fu_1790_p_din1;
    input [63:0] grp_fu_1790_p_dout0;
    output grp_fu_1790_p_ce;
    output [63:0] grp_fu_1794_p_din0;
    output [63:0] grp_fu_1794_p_din1;
    output [4:0] grp_fu_1794_p_opcode;
    input [0:0] grp_fu_1794_p_dout0;
    output grp_fu_1794_p_ce;
    output [63:0] grp_fu_1798_p_din0;
    output [63:0] grp_fu_1798_p_din1;
    input [63:0] grp_fu_1798_p_dout0;
    output grp_fu_1798_p_ce;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg [6:0] p1_address0;
    reg p1_ce0;
    reg [6:0] p1_address1;
    reg p1_ce1;
    reg [5:0] axes1_address0;
    reg axes1_ce0;
    reg [5:0] axes1_address1;
    reg axes1_ce1;
    reg [2:0] p2_0_0_address0;
    reg p2_0_0_ce0;
    reg [2:0] p2_0_1_address0;
    reg p2_0_1_ce0;
    reg [2:0] p2_0_2_address0;
    reg p2_0_2_ce0;
    reg [2:0] p2_1_0_address0;
    reg p2_1_0_ce0;
    reg [2:0] p2_1_1_address0;
    reg p2_1_1_ce0;
    reg [2:0] p2_1_2_address0;
    reg p2_1_2_ce0;
    reg [2:0] p2_2_0_address0;
    reg p2_2_0_ce0;
    reg [2:0] p2_2_1_address0;
    reg p2_2_1_ce0;
    reg [2:0] p2_2_2_address0;
    reg p2_2_2_ce0;
    reg [2:0] p2_3_0_address0;
    reg p2_3_0_ce0;
    reg [2:0] p2_3_1_address0;
    reg p2_3_1_ce0;
    reg [2:0] p2_3_2_address0;
    reg p2_3_2_ce0;
    reg [2:0] p2_4_0_address0;
    reg p2_4_0_ce0;
    reg [2:0] p2_4_1_address0;
    reg p2_4_1_ce0;
    reg [2:0] p2_4_2_address0;
    reg p2_4_2_ce0;
    reg [2:0] p2_5_0_address0;
    reg p2_5_0_ce0;
    reg [2:0] p2_5_1_address0;
    reg p2_5_1_ce0;
    reg [2:0] p2_5_2_address0;
    reg p2_5_2_ce0;
    reg [2:0] p2_6_0_address0;
    reg p2_6_0_ce0;
    reg [2:0] p2_6_1_address0;
    reg p2_6_1_ce0;
    reg [2:0] p2_6_2_address0;
    reg p2_6_2_ce0;
    reg [2:0] p2_7_0_address0;
    reg p2_7_0_ce0;
    reg [2:0] p2_7_1_address0;
    reg p2_7_1_ce0;
    reg [2:0] p2_7_2_address0;
    reg p2_7_2_ce0;
    reg [2:0] p2_8_0_address0;
    reg p2_8_0_ce0;
    reg [2:0] p2_8_1_address0;
    reg p2_8_1_ce0;
    reg [2:0] p2_8_2_address0;
    reg p2_8_2_ce0;
    reg [6:0] axes2_address0;
    reg axes2_ce0;
    reg [6:0] axes2_address1;
    reg axes2_ce1;
    reg [0:0] ap_return;

    (* fsm_encoding = "none" *) reg [103:0] ap_CS_fsm;
    wire ap_CS_fsm_state1;
    reg [63:0] reg_531;
    wire ap_CS_fsm_state3;
    wire ap_CS_fsm_state11;
    reg [63:0] reg_538;
    reg [63:0] reg_545;
    wire ap_CS_fsm_state18;
    wire ap_CS_fsm_state25;
    wire ap_CS_fsm_state32;
    wire ap_CS_fsm_state96;
    reg [63:0] reg_554;
    reg [63:0] reg_562;
    reg [63:0] reg_570;
    reg [63:0] reg_576;
    reg [63:0] reg_582;
    reg [63:0] reg_588;
    wire ap_CS_fsm_state89;
    wire [6:0] mul_ln160_fu_598_p2;
    reg [6:0] mul_ln160_reg_795;
    wire ap_CS_fsm_state2;
    wire [63:0] p2_offset_cast_fu_618_p1;
    reg [63:0] p2_offset_cast_reg_824;
    reg [63:0] y_1_load_reg_860;
    wire ap_CS_fsm_state4;
    reg [63:0] p2_0_1_load_reg_866;
    reg [63:0] y_2_load_reg_872;
    reg [63:0] p1_load_28_reg_877;
    reg [63:0] y_load_reg_882;
    reg [63:0] p2_1_1_load_reg_887;
    wire ap_CS_fsm_state10;
    reg [63:0] p2_0_2_load_reg_912;
    reg [63:0] sub5_i1_reg_918;
    reg [63:0] sub_i2_reg_924;
    reg [63:0] sub5_i2_reg_930;
    reg [63:0] p2_1_2_load_reg_936;
    reg [63:0] mul5_i_i1_reg_941;
    wire [63:0] grp_fu_509_p2;
    reg [63:0] mul_i_i2_reg_946;
    wire [63:0] grp_fu_513_p2;
    reg [63:0] mul5_i_i2_reg_951;
    wire [63:0] grp_fu_526_p2;
    reg [63:0] tmp_6_reg_956;
    wire [0:0] icmp_ln160_fu_702_p2;
    reg [0:0] icmp_ln160_reg_961;
    wire ap_CS_fsm_state97;
    wire [0:0] icmp_ln160_1_fu_708_p2;
    reg [0:0] icmp_ln160_1_reg_966;
    wire [0:0] icmp_ln160_2_fu_714_p2;
    reg [0:0] icmp_ln160_2_reg_971;
    wire [0:0] icmp_ln160_3_fu_720_p2;
    reg [0:0] icmp_ln160_3_reg_976;
    wire [0:0] and_ln160_1_fu_740_p2;
    reg [0:0] and_ln160_1_reg_981;
    wire ap_CS_fsm_state98;
    wire [5:0] sub_ln179_fu_760_p2;
    reg [5:0] sub_ln179_reg_985;
    wire ap_CS_fsm_state99;
    wire [4:0] empty_fu_780_p2;
    reg [4:0] empty_reg_990;
    wire [0:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return;
    reg [0:0] targetBlock_reg_995;
    wire ap_CS_fsm_state100;
    wire [0:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return;
    reg [0:0] targetBlock1_reg_999;
    wire ap_CS_fsm_state102;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_idle;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_ready;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce1;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_ce0;
    wire [5:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce0;
    wire [5:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_idle;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_ready;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce1;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_done;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_idle;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_ready;
    wire   [5:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce0;
    wire   [5:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce1;
    wire   [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce0;
    wire   [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce1;
    wire   [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address0;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce0;
    wire   [6:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address1;
    wire grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce1;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_ce0;
    wire   [2:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_address0;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_ce0;
    wire   [0:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_return;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din1;
    wire   [0:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_opcode;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_ce;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din1;
    wire   [0:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_opcode;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_ce;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_ce;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_ce;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_ce;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din0;
    wire   [63:0] grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din1;
    wire    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_ce;
    reg [0:0] ap_phi_mux_retval_8_phi_fu_259_p8;
    reg [0:0] retval_8_reg_255;
    wire ap_CS_fsm_state104;
    reg ap_predicate_op535_call_state104;
    reg ap_block_state104_on_subcall_done;
    reg grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg;
    reg grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg;
    wire ap_CS_fsm_state101;
    reg    grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg;
    wire ap_CS_fsm_state103;
    wire [63:0] zext_ln160_2_fu_604_p1;
    wire [63:0] zext_ln155_fu_613_p1;
    wire [63:0] zext_ln160_3_fu_631_p1;
    wire [63:0] zext_ln155_2_fu_641_p1;
    wire [63:0] zext_ln155_1_fu_651_p1;
    wire [63:0] zext_ln155_3_fu_661_p1;
    reg [63:0] grp_fu_469_p0;
    reg [63:0] grp_fu_469_p1;
    wire ap_CS_fsm_state5;
    wire ap_CS_fsm_state12;
    wire ap_CS_fsm_state19;
    wire ap_CS_fsm_state26;
    wire ap_CS_fsm_state90;
    reg [63:0] grp_fu_473_p0;
    reg [63:0] grp_fu_473_p1;
    reg [63:0] grp_fu_477_p0;
    reg [63:0] grp_fu_477_p1;
    reg [63:0] grp_fu_493_p0;
    reg [63:0] grp_fu_493_p1;
    reg [63:0] grp_fu_497_p0;
    reg [63:0] grp_fu_497_p1;
    reg [63:0] grp_fu_501_p0;
    reg [63:0] grp_fu_501_p1;
    reg [63:0] grp_fu_505_p0;
    reg [63:0] grp_fu_505_p1;
    reg [63:0] grp_fu_521_p1;
    wire ap_CS_fsm_state33;
    wire ap_CS_fsm_state40;
    wire [1:0] mul_ln160_fu_598_p0;
    wire [5:0] mul_ln160_fu_598_p1;
    wire [6:0] add_ln155_fu_608_p2;
    wire [6:0] add_ln160_fu_626_p2;
    wire [6:0] add_ln155_2_fu_636_p2;
    wire [6:0] add_ln155_1_fu_646_p2;
    wire [6:0] add_ln155_3_fu_656_p2;
    wire [63:0] bitcast_ln160_fu_666_p1;
    wire [63:0] bitcast_ln160_1_fu_684_p1;
    wire [10:0] tmp_304_fu_670_p4;
    wire [51:0] trunc_ln160_fu_680_p1;
    wire [10:0] tmp_305_fu_688_p4;
    wire [51:0] trunc_ln160_1_fu_698_p1;
    wire [0:0] or_ln160_fu_726_p2;
    wire [0:0] or_ln160_1_fu_730_p2;
    wire [0:0] and_ln160_fu_734_p2;
    wire [4:0] tmp_49_fu_749_p3;
    wire [5:0] zext_ln179_4_fu_756_p1;
    wire [5:0] zext_ln179_fu_746_p1;
    wire [3:0] tmp_50_fu_769_p3;
    wire [4:0] tmp_50_cast_fu_776_p1;
    wire [4:0] zext_ln160_fu_766_p1;
    reg [1:0] grp_fu_469_opcode;
    reg grp_fu_469_ce;
    reg [1:0] grp_fu_473_opcode;
    reg grp_fu_473_ce;
    reg [1:0] grp_fu_477_opcode;
    reg grp_fu_493_ce;
    reg grp_fu_497_ce;
    reg grp_fu_501_ce;
    reg grp_fu_505_ce;
    reg [0:0] ap_return_preg;
    reg [103:0] ap_NS_fsm;
    reg ap_ST_fsm_state1_blk;
    wire ap_ST_fsm_state2_blk;
    wire ap_ST_fsm_state3_blk;
    wire ap_ST_fsm_state4_blk;
    wire ap_ST_fsm_state5_blk;
    wire ap_ST_fsm_state6_blk;
    wire ap_ST_fsm_state7_blk;
    wire ap_ST_fsm_state8_blk;
    wire ap_ST_fsm_state9_blk;
    wire ap_ST_fsm_state10_blk;
    wire ap_ST_fsm_state11_blk;
    wire ap_ST_fsm_state12_blk;
    wire ap_ST_fsm_state13_blk;
    wire ap_ST_fsm_state14_blk;
    wire ap_ST_fsm_state15_blk;
    wire ap_ST_fsm_state16_blk;
    wire ap_ST_fsm_state17_blk;
    wire ap_ST_fsm_state18_blk;
    wire ap_ST_fsm_state19_blk;
    wire ap_ST_fsm_state20_blk;
    wire ap_ST_fsm_state21_blk;
    wire ap_ST_fsm_state22_blk;
    wire ap_ST_fsm_state23_blk;
    wire ap_ST_fsm_state24_blk;
    wire ap_ST_fsm_state25_blk;
    wire ap_ST_fsm_state26_blk;
    wire ap_ST_fsm_state27_blk;
    wire ap_ST_fsm_state28_blk;
    wire ap_ST_fsm_state29_blk;
    wire ap_ST_fsm_state30_blk;
    wire ap_ST_fsm_state31_blk;
    wire ap_ST_fsm_state32_blk;
    wire ap_ST_fsm_state33_blk;
    wire ap_ST_fsm_state34_blk;
    wire ap_ST_fsm_state35_blk;
    wire ap_ST_fsm_state36_blk;
    wire ap_ST_fsm_state37_blk;
    wire ap_ST_fsm_state38_blk;
    wire ap_ST_fsm_state39_blk;
    wire ap_ST_fsm_state40_blk;
    wire ap_ST_fsm_state41_blk;
    wire ap_ST_fsm_state42_blk;
    wire ap_ST_fsm_state43_blk;
    wire ap_ST_fsm_state44_blk;
    wire ap_ST_fsm_state45_blk;
    wire ap_ST_fsm_state46_blk;
    wire ap_ST_fsm_state47_blk;
    wire ap_ST_fsm_state48_blk;
    wire ap_ST_fsm_state49_blk;
    wire ap_ST_fsm_state50_blk;
    wire ap_ST_fsm_state51_blk;
    wire ap_ST_fsm_state52_blk;
    wire ap_ST_fsm_state53_blk;
    wire ap_ST_fsm_state54_blk;
    wire ap_ST_fsm_state55_blk;
    wire ap_ST_fsm_state56_blk;
    wire ap_ST_fsm_state57_blk;
    wire ap_ST_fsm_state58_blk;
    wire ap_ST_fsm_state59_blk;
    wire ap_ST_fsm_state60_blk;
    wire ap_ST_fsm_state61_blk;
    wire ap_ST_fsm_state62_blk;
    wire ap_ST_fsm_state63_blk;
    wire ap_ST_fsm_state64_blk;
    wire ap_ST_fsm_state65_blk;
    wire ap_ST_fsm_state66_blk;
    wire ap_ST_fsm_state67_blk;
    wire ap_ST_fsm_state68_blk;
    wire ap_ST_fsm_state69_blk;
    wire ap_ST_fsm_state70_blk;
    wire ap_ST_fsm_state71_blk;
    wire ap_ST_fsm_state72_blk;
    wire ap_ST_fsm_state73_blk;
    wire ap_ST_fsm_state74_blk;
    wire ap_ST_fsm_state75_blk;
    wire ap_ST_fsm_state76_blk;
    wire ap_ST_fsm_state77_blk;
    wire ap_ST_fsm_state78_blk;
    wire ap_ST_fsm_state79_blk;
    wire ap_ST_fsm_state80_blk;
    wire ap_ST_fsm_state81_blk;
    wire ap_ST_fsm_state82_blk;
    wire ap_ST_fsm_state83_blk;
    wire ap_ST_fsm_state84_blk;
    wire ap_ST_fsm_state85_blk;
    wire ap_ST_fsm_state86_blk;
    wire ap_ST_fsm_state87_blk;
    wire ap_ST_fsm_state88_blk;
    wire ap_ST_fsm_state89_blk;
    wire ap_ST_fsm_state90_blk;
    wire ap_ST_fsm_state91_blk;
    wire ap_ST_fsm_state92_blk;
    wire ap_ST_fsm_state93_blk;
    wire ap_ST_fsm_state94_blk;
    wire ap_ST_fsm_state95_blk;
    wire ap_ST_fsm_state96_blk;
    wire ap_ST_fsm_state97_blk;
    wire ap_ST_fsm_state98_blk;
    wire ap_ST_fsm_state99_blk;
    reg ap_ST_fsm_state100_blk;
    wire ap_ST_fsm_state101_blk;
    reg ap_ST_fsm_state102_blk;
    wire ap_ST_fsm_state103_blk;
    reg ap_ST_fsm_state104_blk;
    wire [6:0] mul_ln160_fu_598_p00;
    wire ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 104'd1;
        #0 grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg = 1'b0;
        #0 grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg = 1'b0;
        #0
        grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg = 1'b0;
        #0 ap_return_preg = 1'd0;
    end

    main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1 grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start),
        .ap_done(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done),
        .ap_idle(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_idle),
        .ap_ready(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_ready),
        .p1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address0),
        .p1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce0),
        .p1_q0(p1_q0),
        .p1_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address1),
        .p1_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce1),
        .p1_q1(p1_q1),
        .p1_offset(p1_offset),
        .p2_0_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_address0),
        .p2_0_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_ce0),
        .p2_0_0_q0(p2_0_0_q0),
        .p2_0_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_address0),
        .p2_0_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_ce0),
        .p2_0_1_q0(p2_0_1_q0),
        .p2_0_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_address0),
        .p2_0_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_ce0),
        .p2_0_2_q0(p2_0_2_q0),
        .p2_1_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_address0),
        .p2_1_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_ce0),
        .p2_1_0_q0(p2_1_0_q0),
        .p2_1_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_address0),
        .p2_1_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_ce0),
        .p2_1_1_q0(p2_1_1_q0),
        .p2_1_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_address0),
        .p2_1_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_ce0),
        .p2_1_2_q0(p2_1_2_q0),
        .p2_2_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_address0),
        .p2_2_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_ce0),
        .p2_2_0_q0(p2_2_0_q0),
        .p2_2_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_address0),
        .p2_2_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_ce0),
        .p2_2_1_q0(p2_2_1_q0),
        .p2_2_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_address0),
        .p2_2_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_ce0),
        .p2_2_2_q0(p2_2_2_q0),
        .p2_3_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_address0),
        .p2_3_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_ce0),
        .p2_3_0_q0(p2_3_0_q0),
        .p2_3_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_address0),
        .p2_3_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_ce0),
        .p2_3_1_q0(p2_3_1_q0),
        .p2_3_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_address0),
        .p2_3_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_ce0),
        .p2_3_2_q0(p2_3_2_q0),
        .p2_4_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_address0),
        .p2_4_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_ce0),
        .p2_4_0_q0(p2_4_0_q0),
        .p2_4_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_address0),
        .p2_4_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_ce0),
        .p2_4_1_q0(p2_4_1_q0),
        .p2_4_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_address0),
        .p2_4_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_ce0),
        .p2_4_2_q0(p2_4_2_q0),
        .p2_5_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_address0),
        .p2_5_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_ce0),
        .p2_5_0_q0(p2_5_0_q0),
        .p2_5_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_address0),
        .p2_5_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_ce0),
        .p2_5_1_q0(p2_5_1_q0),
        .p2_5_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_address0),
        .p2_5_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_ce0),
        .p2_5_2_q0(p2_5_2_q0),
        .p2_6_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_address0),
        .p2_6_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_ce0),
        .p2_6_0_q0(p2_6_0_q0),
        .p2_6_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_address0),
        .p2_6_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_ce0),
        .p2_6_1_q0(p2_6_1_q0),
        .p2_6_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_address0),
        .p2_6_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_ce0),
        .p2_6_2_q0(p2_6_2_q0),
        .p2_7_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_address0),
        .p2_7_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_ce0),
        .p2_7_0_q0(p2_7_0_q0),
        .p2_7_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_address0),
        .p2_7_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_ce0),
        .p2_7_1_q0(p2_7_1_q0),
        .p2_7_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_address0),
        .p2_7_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_ce0),
        .p2_7_2_q0(p2_7_2_q0),
        .p2_8_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_address0),
        .p2_8_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_ce0),
        .p2_8_0_q0(p2_8_0_q0),
        .p2_8_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_address0),
        .p2_8_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_ce0),
        .p2_8_1_q0(p2_8_1_q0),
        .p2_8_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_address0),
        .p2_8_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_ce0),
        .p2_8_2_q0(p2_8_2_q0),
        .p2_offset(p2_offset),
        .axes1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address0),
        .axes1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce0),
        .axes1_q0(axes1_q0),
        .axes1_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address1),
        .axes1_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce1),
        .axes1_q1(axes1_q1),
        .ap_return(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return)
    );

    main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2 grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start),
        .ap_done(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done),
        .ap_idle(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_idle),
        .ap_ready(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_ready),
        .p1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address0),
        .p1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce0),
        .p1_q0(p1_q0),
        .p1_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address1),
        .p1_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce1),
        .p1_q1(p1_q1),
        .p1_offset(p1_offset),
        .p2_0_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_address0),
        .p2_0_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_ce0),
        .p2_0_0_q0(p2_0_0_q0),
        .p2_0_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_address0),
        .p2_0_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_ce0),
        .p2_0_1_q0(p2_0_1_q0),
        .p2_0_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_address0),
        .p2_0_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_ce0),
        .p2_0_2_q0(p2_0_2_q0),
        .p2_1_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_address0),
        .p2_1_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_ce0),
        .p2_1_0_q0(p2_1_0_q0),
        .p2_1_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_address0),
        .p2_1_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_ce0),
        .p2_1_1_q0(p2_1_1_q0),
        .p2_1_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_address0),
        .p2_1_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_ce0),
        .p2_1_2_q0(p2_1_2_q0),
        .p2_2_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_address0),
        .p2_2_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_ce0),
        .p2_2_0_q0(p2_2_0_q0),
        .p2_2_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_address0),
        .p2_2_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_ce0),
        .p2_2_1_q0(p2_2_1_q0),
        .p2_2_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_address0),
        .p2_2_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_ce0),
        .p2_2_2_q0(p2_2_2_q0),
        .p2_3_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_address0),
        .p2_3_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_ce0),
        .p2_3_0_q0(p2_3_0_q0),
        .p2_3_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_address0),
        .p2_3_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_ce0),
        .p2_3_1_q0(p2_3_1_q0),
        .p2_3_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_address0),
        .p2_3_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_ce0),
        .p2_3_2_q0(p2_3_2_q0),
        .p2_4_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_address0),
        .p2_4_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_ce0),
        .p2_4_0_q0(p2_4_0_q0),
        .p2_4_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_address0),
        .p2_4_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_ce0),
        .p2_4_1_q0(p2_4_1_q0),
        .p2_4_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_address0),
        .p2_4_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_ce0),
        .p2_4_2_q0(p2_4_2_q0),
        .p2_5_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_address0),
        .p2_5_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_ce0),
        .p2_5_0_q0(p2_5_0_q0),
        .p2_5_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_address0),
        .p2_5_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_ce0),
        .p2_5_1_q0(p2_5_1_q0),
        .p2_5_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_address0),
        .p2_5_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_ce0),
        .p2_5_2_q0(p2_5_2_q0),
        .p2_6_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_address0),
        .p2_6_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_ce0),
        .p2_6_0_q0(p2_6_0_q0),
        .p2_6_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_address0),
        .p2_6_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_ce0),
        .p2_6_1_q0(p2_6_1_q0),
        .p2_6_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_address0),
        .p2_6_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_ce0),
        .p2_6_2_q0(p2_6_2_q0),
        .p2_7_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_address0),
        .p2_7_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_ce0),
        .p2_7_0_q0(p2_7_0_q0),
        .p2_7_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_address0),
        .p2_7_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_ce0),
        .p2_7_1_q0(p2_7_1_q0),
        .p2_7_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_address0),
        .p2_7_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_ce0),
        .p2_7_2_q0(p2_7_2_q0),
        .p2_8_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_address0),
        .p2_8_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_ce0),
        .p2_8_0_q0(p2_8_0_q0),
        .p2_8_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_address0),
        .p2_8_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_ce0),
        .p2_8_1_q0(p2_8_1_q0),
        .p2_8_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_address0),
        .p2_8_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_ce0),
        .p2_8_2_q0(p2_8_2_q0),
        .p2_offset(p2_offset),
        .axes2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address0),
        .axes2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce0),
        .axes2_q0(axes2_q0),
        .axes2_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address1),
        .axes2_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce1),
        .axes2_q1(axes2_q1),
        .ap_return(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return)
    );

    main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4 grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start),
        .ap_done(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_done),
        .ap_idle(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_idle),
        .ap_ready(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_ready),
        .empty(empty_reg_990),
        .axes1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address0),
        .axes1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce0),
        .axes1_q0(axes1_q0),
        .axes1_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address1),
        .axes1_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce1),
        .axes1_q1(axes1_q1),
        .sub_ln179(sub_ln179_reg_985),
        .axes2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address0),
        .axes2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce0),
        .axes2_q0(axes2_q0),
        .axes2_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address1),
        .axes2_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce1),
        .axes2_q1(axes2_q1),
        .p1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address0),
        .p1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce0),
        .p1_q0(p1_q0),
        .p1_address1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address1),
        .p1_ce1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce1),
        .p1_q1(p1_q1),
        .p1_offset(p1_offset),
        .p2_0_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_address0),
        .p2_0_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_ce0),
        .p2_0_0_q0(p2_0_0_q0),
        .p2_0_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_address0),
        .p2_0_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_ce0),
        .p2_0_1_q0(p2_0_1_q0),
        .p2_0_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_address0),
        .p2_0_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_ce0),
        .p2_0_2_q0(p2_0_2_q0),
        .p2_1_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_address0),
        .p2_1_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_ce0),
        .p2_1_0_q0(p2_1_0_q0),
        .p2_1_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_address0),
        .p2_1_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_ce0),
        .p2_1_1_q0(p2_1_1_q0),
        .p2_1_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_address0),
        .p2_1_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_ce0),
        .p2_1_2_q0(p2_1_2_q0),
        .p2_2_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_address0),
        .p2_2_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_ce0),
        .p2_2_0_q0(p2_2_0_q0),
        .p2_2_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_address0),
        .p2_2_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_ce0),
        .p2_2_1_q0(p2_2_1_q0),
        .p2_2_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_address0),
        .p2_2_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_ce0),
        .p2_2_2_q0(p2_2_2_q0),
        .p2_3_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_address0),
        .p2_3_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_ce0),
        .p2_3_0_q0(p2_3_0_q0),
        .p2_3_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_address0),
        .p2_3_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_ce0),
        .p2_3_1_q0(p2_3_1_q0),
        .p2_3_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_address0),
        .p2_3_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_ce0),
        .p2_3_2_q0(p2_3_2_q0),
        .p2_4_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_address0),
        .p2_4_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_ce0),
        .p2_4_0_q0(p2_4_0_q0),
        .p2_4_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_address0),
        .p2_4_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_ce0),
        .p2_4_1_q0(p2_4_1_q0),
        .p2_4_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_address0),
        .p2_4_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_ce0),
        .p2_4_2_q0(p2_4_2_q0),
        .p2_5_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_address0),
        .p2_5_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_ce0),
        .p2_5_0_q0(p2_5_0_q0),
        .p2_5_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_address0),
        .p2_5_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_ce0),
        .p2_5_1_q0(p2_5_1_q0),
        .p2_5_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_address0),
        .p2_5_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_ce0),
        .p2_5_2_q0(p2_5_2_q0),
        .p2_6_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_address0),
        .p2_6_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_ce0),
        .p2_6_0_q0(p2_6_0_q0),
        .p2_6_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_address0),
        .p2_6_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_ce0),
        .p2_6_1_q0(p2_6_1_q0),
        .p2_6_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_address0),
        .p2_6_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_ce0),
        .p2_6_2_q0(p2_6_2_q0),
        .p2_7_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_address0),
        .p2_7_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_ce0),
        .p2_7_0_q0(p2_7_0_q0),
        .p2_7_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_address0),
        .p2_7_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_ce0),
        .p2_7_1_q0(p2_7_1_q0),
        .p2_7_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_address0),
        .p2_7_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_ce0),
        .p2_7_2_q0(p2_7_2_q0),
        .p2_8_0_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_address0),
        .p2_8_0_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_ce0),
        .p2_8_0_q0(p2_8_0_q0),
        .p2_8_1_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_address0),
        .p2_8_1_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_ce0),
        .p2_8_1_q0(p2_8_1_q0),
        .p2_8_2_address0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_address0),
        .p2_8_2_ce0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_ce0),
        .p2_8_2_q0(p2_8_2_q0),
        .p2_offset(p2_offset),
        .ap_return(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_return),
        .grp_fu_469_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din0),
        .grp_fu_469_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din1),
        .grp_fu_469_p_opcode(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_opcode),
        .grp_fu_469_p_dout0(grp_fu_1754_p_dout0),
        .grp_fu_469_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_ce),
        .grp_fu_473_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din0),
        .grp_fu_473_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din1),
        .grp_fu_473_p_opcode(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_opcode),
        .grp_fu_473_p_dout0(grp_fu_1762_p_dout0),
        .grp_fu_473_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_ce),
        .grp_fu_493_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din0),
        .grp_fu_493_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din1),
        .grp_fu_493_p_dout0(grp_fu_1758_p_dout0),
        .grp_fu_493_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_ce),
        .grp_fu_497_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din0),
        .grp_fu_497_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din1),
        .grp_fu_497_p_dout0(grp_fu_1782_p_dout0),
        .grp_fu_497_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_ce),
        .grp_fu_501_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din0),
        .grp_fu_501_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din1),
        .grp_fu_501_p_dout0(grp_fu_1786_p_dout0),
        .grp_fu_501_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_ce),
        .grp_fu_505_p_din0(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din0),
        .grp_fu_505_p_din1(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din1),
        .grp_fu_505_p_dout0(grp_fu_1790_p_dout0),
        .grp_fu_505_p_ce(grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_ce)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U1341 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(sub_i2_reg_924),
        .din1(sub_i2_reg_924),
        .ce(1'b1),
        .dout(grp_fu_509_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_x_U1342 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(sub5_i2_reg_930),
        .din1(sub5_i2_reg_930),
        .ce(1'b1),
        .dout(grp_fu_513_p2)
    );

    main_dsqrt_64ns_64ns_64_57_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(57),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsqrt_64ns_64ns_64_57_no_dsp_1_U1345 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd0),
        .din1(reg_562),
        .ce(1'b1),
        .dout(grp_fu_526_p2)
    );

    main_mul_2ns_6ns_7_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(2),
        .din1_WIDTH(6),
        .dout_WIDTH(7)
    ) mul_2ns_6ns_7_1_1_U1346 (
        .din0(mul_ln160_fu_598_p0),
        .din1(mul_ln160_fu_598_p1),
        .dout(mul_ln160_fu_598_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg <= 1'd0;
        end else begin
            if (((1'b0 == ap_block_state104_on_subcall_done) & (1'b1 == ap_CS_fsm_state104))) begin
                ap_return_preg <= ap_phi_mux_retval_8_phi_fu_259_p8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd0 == and_ln160_1_reg_981) & (1'b1 == ap_CS_fsm_state99))) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg <= 1'b1;
            end else if ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_ready == 1'b1)) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state101)) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg <= 1'b1;
            end else if ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_ready == 1'b1)) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state103)) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg <= 1'b1;
            end else if ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_ready == 1'b1)) begin
                grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state100)) | ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state102)) | ((1'd1 == and_ln160_1_reg_981) & (1'b1 == ap_CS_fsm_state99)))) begin
            retval_8_reg_255 <= 1'd0;
        end else if (((1'b0 == ap_block_state104_on_subcall_done) & (1'd0 == and_ln160_1_reg_981) & (targetBlock1_reg_999 == 1'd1) & (targetBlock_reg_995 == 1'd1) & (1'b1 == ap_CS_fsm_state104))) begin
            retval_8_reg_255 <= grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state98)) begin
            and_ln160_1_reg_981 <= and_ln160_1_fu_740_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state99)) begin
            empty_reg_990 <= empty_fu_780_p2;
            sub_ln179_reg_985 <= sub_ln179_fu_760_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state97)) begin
            icmp_ln160_1_reg_966 <= icmp_ln160_1_fu_708_p2;
            icmp_ln160_2_reg_971 <= icmp_ln160_2_fu_714_p2;
            icmp_ln160_3_reg_976 <= icmp_ln160_3_fu_720_p2;
            icmp_ln160_reg_961   <= icmp_ln160_fu_702_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state18)) begin
            mul5_i_i1_reg_941 <= grp_fu_1790_p_dout0;
            mul5_i_i2_reg_951 <= grp_fu_513_p2;
            mul_i_i2_reg_946  <= grp_fu_509_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            mul_ln160_reg_795 <= mul_ln160_fu_598_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            p1_load_28_reg_877 <= p1_q0;
            p2_0_1_load_reg_866 <= p2_0_1_q0;
            p2_1_1_load_reg_887 <= p2_1_1_q0;
            y_1_load_reg_860 <= p2_0_0_q0;
            y_2_load_reg_872 <= p1_q1;
            y_load_reg_882 <= p2_1_0_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            p2_0_2_load_reg_912 <= p2_0_2_q0;
            p2_1_2_load_reg_936 <= p2_1_2_q0;
            sub5_i1_reg_918 <= grp_fu_1770_p_dout0;
            sub5_i2_reg_930 <= grp_fu_1778_p_dout0;
            sub_i2_reg_924 <= grp_fu_1774_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_offset_cast_reg_824[2 : 0] <= p2_offset_cast_fu_618_p1[2 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state3))) begin
            reg_531 <= p1_q1;
            reg_538 <= p1_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state96) | (1'b1 == ap_CS_fsm_state32) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state11))) begin
            reg_545 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state32) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state11))) begin
            reg_554 <= grp_fu_1762_p_dout0;
            reg_562 <= grp_fu_1766_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state18))) begin
            reg_570 <= grp_fu_1758_p_dout0;
            reg_576 <= grp_fu_1782_p_dout0;
            reg_582 <= grp_fu_1786_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state89) | (1'b1 == ap_CS_fsm_state96))) begin
            reg_588 <= grp_fu_1798_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state102)) begin
            targetBlock1_reg_999 <= grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state100)) begin
            targetBlock_reg_995 <= grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state89)) begin
            tmp_6_reg_956 <= grp_fu_526_p2;
        end
    end

    always @(*) begin
        if ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done == 1'b0)) begin
            ap_ST_fsm_state100_blk = 1'b1;
        end else begin
            ap_ST_fsm_state100_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state101_blk = 1'b0;

    always @(*) begin
        if ((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done == 1'b0)) begin
            ap_ST_fsm_state102_blk = 1'b1;
        end else begin
            ap_ST_fsm_state102_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state103_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state104_on_subcall_done)) begin
            ap_ST_fsm_state104_blk = 1'b1;
        end else begin
            ap_ST_fsm_state104_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    assign ap_ST_fsm_state73_blk = 1'b0;

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state75_blk = 1'b0;

    assign ap_ST_fsm_state76_blk = 1'b0;

    assign ap_ST_fsm_state77_blk = 1'b0;

    assign ap_ST_fsm_state78_blk = 1'b0;

    assign ap_ST_fsm_state79_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state80_blk = 1'b0;

    assign ap_ST_fsm_state81_blk = 1'b0;

    assign ap_ST_fsm_state82_blk = 1'b0;

    assign ap_ST_fsm_state83_blk = 1'b0;

    assign ap_ST_fsm_state84_blk = 1'b0;

    assign ap_ST_fsm_state85_blk = 1'b0;

    assign ap_ST_fsm_state86_blk = 1'b0;

    assign ap_ST_fsm_state87_blk = 1'b0;

    assign ap_ST_fsm_state88_blk = 1'b0;

    assign ap_ST_fsm_state89_blk = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state90_blk = 1'b0;

    assign ap_ST_fsm_state91_blk = 1'b0;

    assign ap_ST_fsm_state92_blk = 1'b0;

    assign ap_ST_fsm_state93_blk = 1'b0;

    assign ap_ST_fsm_state94_blk = 1'b0;

    assign ap_ST_fsm_state95_blk = 1'b0;

    assign ap_ST_fsm_state96_blk = 1'b0;

    assign ap_ST_fsm_state97_blk = 1'b0;

    assign ap_ST_fsm_state98_blk = 1'b0;

    assign ap_ST_fsm_state99_blk = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if ((((1'b0 == ap_block_state104_on_subcall_done) & (1'b1 == ap_CS_fsm_state104)) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'd0 == and_ln160_1_reg_981) & (targetBlock1_reg_999 == 1'd1) & (targetBlock_reg_995 == 1'd1) & (1'b1 == ap_CS_fsm_state104))) begin
            ap_phi_mux_retval_8_phi_fu_259_p8 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_return;
        end else begin
            ap_phi_mux_retval_8_phi_fu_259_p8 = retval_8_reg_255;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_state104_on_subcall_done) & (1'b1 == ap_CS_fsm_state104))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_state104_on_subcall_done) & (1'b1 == ap_CS_fsm_state104))) begin
            ap_return = ap_phi_mux_retval_8_phi_fu_259_p8;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            axes1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address0;
        end else begin
            axes1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes1_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_address1;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            axes1_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_address1;
        end else begin
            axes1_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            axes1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce0;
        end else begin
            axes1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes1_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes1_ce1;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            axes1_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_axes1_ce1;
        end else begin
            axes1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            axes2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address0;
        end else begin
            axes2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes2_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_address1;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            axes2_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_address1;
        end else begin
            axes2_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            axes2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce0;
        end else begin
            axes2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            axes2_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_axes2_ce1;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            axes2_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_axes2_ce1;
        end else begin
            axes2_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_469_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_ce;
        end else begin
            grp_fu_469_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_469_opcode = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_opcode;
        end else if (((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5))) begin
            grp_fu_469_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state90) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state19))) begin
            grp_fu_469_opcode = 2'd0;
        end else begin
            grp_fu_469_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_469_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state90)) begin
            grp_fu_469_p0 = reg_588;
        end else if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_469_p0 = reg_545;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_469_p0 = reg_570;
        end else if (((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5))) begin
            grp_fu_469_p0 = reg_531;
        end else begin
            grp_fu_469_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_469_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_469_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state90)) begin
            grp_fu_469_p1 = tmp_6_reg_956;
        end else if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_469_p1 = reg_570;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_469_p1 = reg_576;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_469_p1 = p2_0_2_load_reg_912;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_469_p1 = y_1_load_reg_860;
        end else begin
            grp_fu_469_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_473_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_ce;
        end else begin
            grp_fu_473_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_473_opcode = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_opcode;
        end else if (((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5))) begin
            grp_fu_473_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state19))) begin
            grp_fu_473_opcode = 2'd0;
        end else begin
            grp_fu_473_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_473_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_473_p0 = reg_554;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_473_p0 = reg_582;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_473_p0 = reg_531;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_473_p0 = reg_538;
        end else begin
            grp_fu_473_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_473_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_473_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_473_p1 = reg_576;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_473_p1 = mul5_i_i1_reg_941;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_473_p1 = reg_538;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_473_p1 = p2_0_1_load_reg_866;
        end else begin
            grp_fu_473_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5))) begin
            grp_fu_477_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state19))) begin
            grp_fu_477_opcode = 2'd0;
        end else begin
            grp_fu_477_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_477_p0 = reg_562;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_477_p0 = mul_i_i2_reg_946;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_477_p0 = p2_0_2_load_reg_912;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_477_p0 = reg_531;
        end else begin
            grp_fu_477_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state26)) begin
            grp_fu_477_p1 = reg_582;
        end else if ((1'b1 == ap_CS_fsm_state19)) begin
            grp_fu_477_p1 = mul5_i_i2_reg_951;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_477_p1 = p2_1_2_load_reg_936;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_477_p1 = y_2_load_reg_872;
        end else begin
            grp_fu_477_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_493_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_ce;
        end else begin
            grp_fu_493_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_493_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din0;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_493_p0 = reg_545;
        end else begin
            grp_fu_493_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_493_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_493_p_din1;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_493_p1 = reg_545;
        end else begin
            grp_fu_493_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_497_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_ce;
        end else begin
            grp_fu_497_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_497_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din0;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_497_p0 = reg_554;
        end else begin
            grp_fu_497_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_497_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_497_p_din1;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_497_p1 = reg_554;
        end else begin
            grp_fu_497_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_501_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_ce;
        end else begin
            grp_fu_501_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_501_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din0;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_501_p0 = reg_562;
        end else begin
            grp_fu_501_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_501_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_501_p_din1;
        end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state12))) begin
            grp_fu_501_p1 = reg_562;
        end else begin
            grp_fu_501_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_505_ce = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_ce;
        end else begin
            grp_fu_505_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_505_p0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_505_p0 = sub5_i1_reg_918;
        end else begin
            grp_fu_505_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state104)) begin
            grp_fu_505_p1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_grp_fu_505_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_505_p1 = sub5_i1_reg_918;
        end else begin
            grp_fu_505_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state40)) begin
            grp_fu_521_p1 = reg_545;
        end else if ((1'b1 == ap_CS_fsm_state33)) begin
            grp_fu_521_p1 = reg_554;
        end else begin
            grp_fu_521_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p1_address0 = zext_ln155_3_fu_661_p1;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            p1_address0 = zext_ln155_2_fu_641_p1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            p1_address0 = zext_ln155_fu_613_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address0;
        end else begin
            p1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p1_address1 = zext_ln155_1_fu_651_p1;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            p1_address1 = zext_ln160_3_fu_631_p1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            p1_address1 = zext_ln160_2_fu_604_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p1_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_address1;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p1_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_address1;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p1_address1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_address1;
        end else begin
            p1_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3))) begin
            p1_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce0;
        end else begin
            p1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3))) begin
            p1_ce1 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p1_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p1_ce1;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p1_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p1_ce1;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p1_ce1 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p1_ce1;
        end else begin
            p1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_0_0_address0 = p2_offset_cast_fu_618_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_address0;
        end else begin
            p2_0_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_0_0_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_0_ce0;
        end else begin
            p2_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_0_1_address0 = p2_offset_cast_fu_618_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_address0;
        end else begin
            p2_0_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_0_1_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_1_ce0;
        end else begin
            p2_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p2_0_2_address0 = p2_offset_cast_reg_824;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_address0;
        end else begin
            p2_0_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p2_0_2_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_0_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_0_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_0_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_0_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_0_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_0_2_ce0;
        end else begin
            p2_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_1_0_address0 = p2_offset_cast_fu_618_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_address0;
        end else begin
            p2_1_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_1_0_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_0_ce0;
        end else begin
            p2_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_1_1_address0 = p2_offset_cast_fu_618_p1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_address0;
        end else begin
            p2_1_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            p2_1_1_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_1_ce0;
        end else begin
            p2_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p2_1_2_address0 = p2_offset_cast_reg_824;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_address0;
        end else begin
            p2_1_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            p2_1_2_ce0 = 1'b1;
        end else if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_1_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_1_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_1_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_1_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_1_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_1_2_ce0;
        end else begin
            p2_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_address0;
        end else begin
            p2_2_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_0_ce0;
        end else begin
            p2_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_address0;
        end else begin
            p2_2_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_1_ce0;
        end else begin
            p2_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_address0;
        end else begin
            p2_2_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_2_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_2_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_2_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_2_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_2_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_2_2_ce0;
        end else begin
            p2_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_address0;
        end else begin
            p2_3_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_0_ce0;
        end else begin
            p2_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_address0;
        end else begin
            p2_3_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_1_ce0;
        end else begin
            p2_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_address0;
        end else begin
            p2_3_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_3_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_3_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_3_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_3_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_3_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_3_2_ce0;
        end else begin
            p2_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_address0;
        end else begin
            p2_4_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_0_ce0;
        end else begin
            p2_4_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_address0;
        end else begin
            p2_4_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_1_ce0;
        end else begin
            p2_4_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_address0;
        end else begin
            p2_4_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_4_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_4_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_4_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_4_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_4_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_4_2_ce0;
        end else begin
            p2_4_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_address0;
        end else begin
            p2_5_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_0_ce0;
        end else begin
            p2_5_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_address0;
        end else begin
            p2_5_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_1_ce0;
        end else begin
            p2_5_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_address0;
        end else begin
            p2_5_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_5_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_5_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_5_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_5_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_5_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_5_2_ce0;
        end else begin
            p2_5_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_address0;
        end else begin
            p2_6_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_0_ce0;
        end else begin
            p2_6_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_address0;
        end else begin
            p2_6_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_1_ce0;
        end else begin
            p2_6_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_address0;
        end else begin
            p2_6_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_6_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_6_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_6_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_6_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_6_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_6_2_ce0;
        end else begin
            p2_6_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_address0;
        end else begin
            p2_7_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_0_ce0;
        end else begin
            p2_7_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_address0;
        end else begin
            p2_7_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_1_ce0;
        end else begin
            p2_7_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_address0;
        end else begin
            p2_7_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_7_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_7_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_7_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_7_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_7_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_7_2_ce0;
        end else begin
            p2_7_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_0_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_address0;
        end else begin
            p2_8_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_0_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_0_ce0;
        end else begin
            p2_8_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_1_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_address0;
        end else begin
            p2_8_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_1_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_1_ce0;
        end else begin
            p2_8_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_2_address0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_address0;
        end else begin
            p2_8_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_predicate_op535_call_state104 == 1'b1) & (1'b1 == ap_CS_fsm_state104))) begin
            p2_8_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_p2_8_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state102)) begin
            p2_8_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_p2_8_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            p2_8_2_ce0 = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_p2_8_2_ce0;
        end else begin
            p2_8_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end
            ap_ST_fsm_state78: begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
            ap_ST_fsm_state79: begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end
            ap_ST_fsm_state80: begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
            ap_ST_fsm_state81: begin
                ap_NS_fsm = ap_ST_fsm_state82;
            end
            ap_ST_fsm_state82: begin
                ap_NS_fsm = ap_ST_fsm_state83;
            end
            ap_ST_fsm_state83: begin
                ap_NS_fsm = ap_ST_fsm_state84;
            end
            ap_ST_fsm_state84: begin
                ap_NS_fsm = ap_ST_fsm_state85;
            end
            ap_ST_fsm_state85: begin
                ap_NS_fsm = ap_ST_fsm_state86;
            end
            ap_ST_fsm_state86: begin
                ap_NS_fsm = ap_ST_fsm_state87;
            end
            ap_ST_fsm_state87: begin
                ap_NS_fsm = ap_ST_fsm_state88;
            end
            ap_ST_fsm_state88: begin
                ap_NS_fsm = ap_ST_fsm_state89;
            end
            ap_ST_fsm_state89: begin
                ap_NS_fsm = ap_ST_fsm_state90;
            end
            ap_ST_fsm_state90: begin
                ap_NS_fsm = ap_ST_fsm_state91;
            end
            ap_ST_fsm_state91: begin
                ap_NS_fsm = ap_ST_fsm_state92;
            end
            ap_ST_fsm_state92: begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end
            ap_ST_fsm_state93: begin
                ap_NS_fsm = ap_ST_fsm_state94;
            end
            ap_ST_fsm_state94: begin
                ap_NS_fsm = ap_ST_fsm_state95;
            end
            ap_ST_fsm_state95: begin
                ap_NS_fsm = ap_ST_fsm_state96;
            end
            ap_ST_fsm_state96: begin
                ap_NS_fsm = ap_ST_fsm_state97;
            end
            ap_ST_fsm_state97: begin
                ap_NS_fsm = ap_ST_fsm_state98;
            end
            ap_ST_fsm_state98: begin
                ap_NS_fsm = ap_ST_fsm_state99;
            end
            ap_ST_fsm_state99: begin
                if (((1'd1 == and_ln160_1_reg_981) & (1'b1 == ap_CS_fsm_state99))) begin
                    ap_NS_fsm = ap_ST_fsm_state104;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state100;
                end
            end
            ap_ST_fsm_state100: begin
                if (((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state100))) begin
                    ap_NS_fsm = ap_ST_fsm_state104;
                end else if (((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_return == 1'd1) & (1'b1 == ap_CS_fsm_state100))) begin
                    ap_NS_fsm = ap_ST_fsm_state101;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state100;
                end
            end
            ap_ST_fsm_state101: begin
                ap_NS_fsm = ap_ST_fsm_state102;
            end
            ap_ST_fsm_state102: begin
                if (((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state102))) begin
                    ap_NS_fsm = ap_ST_fsm_state104;
                end else if (((grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_done == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_return == 1'd1) & (1'b1 == ap_CS_fsm_state102))) begin
                    ap_NS_fsm = ap_ST_fsm_state103;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state102;
                end
            end
            ap_ST_fsm_state103: begin
                ap_NS_fsm = ap_ST_fsm_state104;
            end
            ap_ST_fsm_state104: begin
                if (((1'b0 == ap_block_state104_on_subcall_done) & (1'b1 == ap_CS_fsm_state104))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state104;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln155_1_fu_646_p2 = (mul_ln160_reg_795 + 7'd2);

    assign add_ln155_2_fu_636_p2 = (mul_ln160_reg_795 + 7'd4);

    assign add_ln155_3_fu_656_p2 = (mul_ln160_reg_795 + 7'd5);

    assign add_ln155_fu_608_p2 = (mul_ln160_reg_795 + 7'd1);

    assign add_ln160_fu_626_p2 = (mul_ln160_reg_795 + 7'd3);

    assign and_ln160_1_fu_740_p2 = (grp_fu_1794_p_dout0 & and_ln160_fu_734_p2);

    assign and_ln160_fu_734_p2 = (or_ln160_fu_726_p2 & or_ln160_1_fu_730_p2);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state100 = ap_CS_fsm[32'd99];

    assign ap_CS_fsm_state101 = ap_CS_fsm[32'd100];

    assign ap_CS_fsm_state102 = ap_CS_fsm[32'd101];

    assign ap_CS_fsm_state103 = ap_CS_fsm[32'd102];

    assign ap_CS_fsm_state104 = ap_CS_fsm[32'd103];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state40 = ap_CS_fsm[32'd39];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state89 = ap_CS_fsm[32'd88];

    assign ap_CS_fsm_state90 = ap_CS_fsm[32'd89];

    assign ap_CS_fsm_state96 = ap_CS_fsm[32'd95];

    assign ap_CS_fsm_state97 = ap_CS_fsm[32'd96];

    assign ap_CS_fsm_state98 = ap_CS_fsm[32'd97];

    assign ap_CS_fsm_state99 = ap_CS_fsm[32'd98];

    always @(*) begin
        ap_block_state104_on_subcall_done = ((ap_predicate_op535_call_state104 == 1'b1) & (grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_done == 1'b0));
    end

    always @(*) begin
        ap_predicate_op535_call_state104 = ((1'd0 == and_ln160_1_reg_981) & (targetBlock1_reg_999 == 1'd1) & (targetBlock_reg_995 == 1'd1));
    end

    assign bitcast_ln160_1_fu_684_p1 = reg_545;

    assign bitcast_ln160_fu_666_p1 = reg_588;

    assign empty_fu_780_p2 = (tmp_50_cast_fu_776_p1 - zext_ln160_fu_766_p1);

    assign grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1_fu_272_ap_start_reg;

    assign grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_171_2_fu_336_ap_start_reg;

    assign grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start = grp_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4_fu_400_ap_start_reg;

    assign grp_fu_1754_p_ce = grp_fu_469_ce;

    assign grp_fu_1754_p_din0 = grp_fu_469_p0;

    assign grp_fu_1754_p_din1 = grp_fu_469_p1;

    assign grp_fu_1754_p_opcode = grp_fu_469_opcode;

    assign grp_fu_1758_p_ce = grp_fu_493_ce;

    assign grp_fu_1758_p_din0 = grp_fu_493_p0;

    assign grp_fu_1758_p_din1 = grp_fu_493_p1;

    assign grp_fu_1762_p_ce = grp_fu_473_ce;

    assign grp_fu_1762_p_din0 = grp_fu_473_p0;

    assign grp_fu_1762_p_din1 = grp_fu_473_p1;

    assign grp_fu_1762_p_opcode = grp_fu_473_opcode;

    assign grp_fu_1766_p_ce = 1'b1;

    assign grp_fu_1766_p_din0 = grp_fu_477_p0;

    assign grp_fu_1766_p_din1 = grp_fu_477_p1;

    assign grp_fu_1766_p_opcode = grp_fu_477_opcode;

    assign grp_fu_1770_p_ce = 1'b1;

    assign grp_fu_1770_p_din0 = reg_538;

    assign grp_fu_1770_p_din1 = p1_load_28_reg_877;

    assign grp_fu_1770_p_opcode = 2'd1;

    assign grp_fu_1774_p_ce = 1'b1;

    assign grp_fu_1774_p_din0 = y_1_load_reg_860;

    assign grp_fu_1774_p_din1 = y_load_reg_882;

    assign grp_fu_1774_p_opcode = 2'd1;

    assign grp_fu_1778_p_ce = 1'b1;

    assign grp_fu_1778_p_din0 = p2_0_1_load_reg_866;

    assign grp_fu_1778_p_din1 = p2_1_1_load_reg_887;

    assign grp_fu_1778_p_opcode = 2'd1;

    assign grp_fu_1782_p_ce = grp_fu_497_ce;

    assign grp_fu_1782_p_din0 = grp_fu_497_p0;

    assign grp_fu_1782_p_din1 = grp_fu_497_p1;

    assign grp_fu_1786_p_ce = grp_fu_501_ce;

    assign grp_fu_1786_p_din0 = grp_fu_501_p0;

    assign grp_fu_1786_p_din1 = grp_fu_501_p1;

    assign grp_fu_1790_p_ce = grp_fu_505_ce;

    assign grp_fu_1790_p_din0 = grp_fu_505_p0;

    assign grp_fu_1790_p_din1 = grp_fu_505_p1;

    assign grp_fu_1794_p_ce = 1'b1;

    assign grp_fu_1794_p_din0 = reg_588;

    assign grp_fu_1794_p_din1 = reg_545;

    assign grp_fu_1794_p_opcode = 5'd2;

    assign grp_fu_1798_p_ce = 1'b1;

    assign grp_fu_1798_p_din0 = 64'd0;

    assign grp_fu_1798_p_din1 = grp_fu_521_p1;

    assign icmp_ln160_1_fu_708_p2 = ((trunc_ln160_fu_680_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln160_2_fu_714_p2 = ((tmp_305_fu_688_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln160_3_fu_720_p2 = ((trunc_ln160_1_fu_698_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln160_fu_702_p2 = ((tmp_304_fu_670_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign mul_ln160_fu_598_p0 = mul_ln160_fu_598_p00;

    assign mul_ln160_fu_598_p00 = p1_offset;

    assign mul_ln160_fu_598_p1 = 7'd27;

    assign or_ln160_1_fu_730_p2 = (icmp_ln160_3_reg_976 | icmp_ln160_2_reg_971);

    assign or_ln160_fu_726_p2 = (icmp_ln160_reg_961 | icmp_ln160_1_reg_966);

    assign p2_offset_cast_fu_618_p1 = p2_offset;

    assign sub_ln179_fu_760_p2 = (zext_ln179_4_fu_756_p1 - zext_ln179_fu_746_p1);

    assign tmp_304_fu_670_p4 = {{bitcast_ln160_fu_666_p1[62:52]}};

    assign tmp_305_fu_688_p4 = {{bitcast_ln160_1_fu_684_p1[62:52]}};

    assign tmp_49_fu_749_p3 = {{p2_offset}, {2'd0}};

    assign tmp_50_cast_fu_776_p1 = tmp_50_fu_769_p3;

    assign tmp_50_fu_769_p3 = {{p1_offset}, {2'd0}};

    assign trunc_ln160_1_fu_698_p1 = bitcast_ln160_1_fu_684_p1[51:0];

    assign trunc_ln160_fu_680_p1 = bitcast_ln160_fu_666_p1[51:0];

    assign zext_ln155_1_fu_651_p1 = add_ln155_1_fu_646_p2;

    assign zext_ln155_2_fu_641_p1 = add_ln155_2_fu_636_p2;

    assign zext_ln155_3_fu_661_p1 = add_ln155_3_fu_656_p2;

    assign zext_ln155_fu_613_p1 = add_ln155_fu_608_p2;

    assign zext_ln160_2_fu_604_p1 = mul_ln160_reg_795;

    assign zext_ln160_3_fu_631_p1 = add_ln160_fu_626_p2;

    assign zext_ln160_fu_766_p1 = p1_offset;

    assign zext_ln179_4_fu_756_p1 = tmp_49_fu_749_p3;

    assign zext_ln179_fu_746_p1 = p2_offset;

    always @(posedge ap_clk) begin
        p2_offset_cast_reg_824[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_cuboidCuboidCollision_double_s
