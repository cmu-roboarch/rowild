/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_rpyxyzToH_double_2 (
    ap_clk,
    ap_rst,
    x,
    ap_return_0,
    ap_return_1,
    ap_return_2,
    ap_return_3,
    ap_return_4,
    ap_return_5,
    ap_return_6,
    ap_return_7,
    ap_return_8,
    ap_return_9,
    ap_return_10,
    ap_return_11
);


    input ap_clk;
    input ap_rst;
    input [63:0] x;
    output [63:0] ap_return_0;
    output [63:0] ap_return_1;
    output [63:0] ap_return_2;
    output [63:0] ap_return_3;
    output [63:0] ap_return_4;
    output [63:0] ap_return_5;
    output [63:0] ap_return_6;
    output [63:0] ap_return_7;
    output [63:0] ap_return_8;
    output [63:0] ap_return_9;
    output [63:0] ap_return_10;
    output [63:0] ap_return_11;

    reg   [63:0] x_read_reg_532;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] x_read_reg_532_pp0_iter1_reg;
    reg   [63:0] x_read_reg_532_pp0_iter2_reg;
    reg   [63:0] x_read_reg_532_pp0_iter3_reg;
    reg   [63:0] x_read_reg_532_pp0_iter4_reg;
    reg   [63:0] x_read_reg_532_pp0_iter5_reg;
    reg   [63:0] x_read_reg_532_pp0_iter6_reg;
    reg   [63:0] x_read_reg_532_pp0_iter7_reg;
    reg   [63:0] x_read_reg_532_pp0_iter8_reg;
    reg   [63:0] x_read_reg_532_pp0_iter9_reg;
    reg   [63:0] x_read_reg_532_pp0_iter10_reg;
    reg   [63:0] x_read_reg_532_pp0_iter11_reg;
    reg   [63:0] x_read_reg_532_pp0_iter12_reg;
    reg   [63:0] x_read_reg_532_pp0_iter13_reg;
    reg   [63:0] x_read_reg_532_pp0_iter14_reg;
    reg   [63:0] x_read_reg_532_pp0_iter15_reg;
    reg   [63:0] x_read_reg_532_pp0_iter16_reg;
    reg   [63:0] x_read_reg_532_pp0_iter17_reg;
    reg   [63:0] x_read_reg_532_pp0_iter18_reg;
    reg   [63:0] x_read_reg_532_pp0_iter19_reg;
    reg   [63:0] x_read_reg_532_pp0_iter20_reg;
    wire   [63:0] grp_fu_354_p2;
    reg   [63:0] mul_i_0_0_3_reg_538;
    wire   [63:0] grp_fu_18_p2;
    reg   [63:0] add_i_0_0_3_reg_544;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter14_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter15_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter16_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter17_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter18_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter19_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter20_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter21_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter22_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter23_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter24_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter25_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter26_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter27_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter28_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter29_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter30_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter31_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter32_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter33_reg;
    reg   [63:0] add_i_0_0_3_reg_544_pp0_iter34_reg;
    wire   [63:0] grp_fu_23_p2;
    reg   [63:0] add_i_0_1_3_reg_553;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter14_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter15_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter16_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter17_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter18_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter19_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter20_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter21_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter22_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter23_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter24_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter25_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter26_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter27_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter28_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter29_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter30_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter31_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter32_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter33_reg;
    reg   [63:0] add_i_0_1_3_reg_553_pp0_iter34_reg;
    wire   [63:0] grp_fu_28_p2;
    reg   [63:0] add_i1_reg_565;
    wire   [63:0] grp_fu_360_p2;
    reg   [63:0] mul_i1_0_0_1_reg_570;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter21_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter22_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter23_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter24_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter25_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter26_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter27_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter28_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter29_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter30_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter31_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter32_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter33_reg;
    reg   [63:0] mul_i1_0_0_1_reg_570_pp0_iter34_reg;
    wire   [63:0] grp_fu_365_p2;
    reg   [63:0] mul_i1_0_1_reg_583;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter21_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter22_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter23_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter24_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter25_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter26_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter27_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter28_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter29_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter30_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter31_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter32_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter33_reg;
    reg   [63:0] mul_i1_0_1_reg_583_pp0_iter34_reg;
    wire   [63:0] grp_fu_33_p2;
    reg   [63:0] add_i_0_3_3_reg_592;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter28_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter29_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter30_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter31_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter32_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter33_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter34_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter35_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter36_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter37_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter38_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter39_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter40_reg;
    reg   [63:0] add_i_0_3_3_reg_592_pp0_iter41_reg;
    wire   [63:0] grp_fu_38_p2;
    reg   [63:0] add_i1_0_0_1_reg_600;
    wire   [63:0] grp_fu_370_p2;
    reg   [63:0] mul_i1_0_0_2_reg_605;
    wire   [63:0] grp_fu_42_p2;
    reg   [63:0] add_i1_0_1_reg_611;
    wire   [63:0] grp_fu_47_p2;
    reg   [63:0] add_i1_1_0_1_reg_617;
    wire   [63:0] grp_fu_51_p2;
    reg   [63:0] add_i1_1_1_reg_622;
    wire   [63:0] grp_fu_56_p2;
    reg   [63:0] add_i1_2_0_1_reg_630;
    wire   [63:0] grp_fu_375_p2;
    reg   [63:0] mul_i1_2_0_2_reg_635;
    wire   [63:0] grp_fu_60_p2;
    reg   [63:0] add_i1_0_0_2_reg_640;
    wire   [63:0] grp_fu_380_p2;
    reg   [63:0] mul_i1_0_0_3_reg_645;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter35_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter36_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter37_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter38_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter39_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter40_reg;
    reg   [63:0] mul_i1_0_0_3_reg_645_pp0_iter41_reg;
    wire   [63:0] grp_fu_64_p2;
    reg   [63:0] add_i1_0_1_1_reg_658;
    wire   [63:0] grp_fu_68_p2;
    reg   [63:0] add_i1_0_2_1_reg_663;
    wire   [63:0] grp_fu_72_p2;
    reg   [63:0] add_i1_1_0_2_reg_669;
    wire   [63:0] grp_fu_76_p2;
    reg   [63:0] add_i1_1_1_1_reg_674;
    wire   [63:0] grp_fu_80_p2;
    reg   [63:0] add_i1_1_2_1_reg_679;
    wire   [63:0] grp_fu_84_p2;
    reg   [63:0] add_i1_2_0_2_reg_685;
    wire   [63:0] grp_fu_88_p2;
    reg   [63:0] add_i1_2_1_1_reg_690;
    wire   [63:0] grp_fu_92_p2;
    reg   [63:0] add_i1_2_2_1_reg_695;
    wire   [63:0] grp_fu_96_p2;
    reg   [63:0] add_i1_0_0_3_reg_701;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter42_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter43_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter44_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter45_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter46_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter47_reg;
    reg   [63:0] add_i1_0_0_3_reg_701_pp0_iter48_reg;
    wire   [63:0] grp_fu_100_p2;
    reg   [63:0] add_i1_0_1_2_reg_707;
    wire   [63:0] grp_fu_104_p2;
    reg   [63:0] add_i1_0_2_2_reg_712;
    wire   [63:0] grp_fu_108_p2;
    reg   [63:0] add_i1_0_3_2_reg_717;
    wire   [63:0] grp_fu_112_p2;
    reg   [63:0] add_i1_1_0_3_reg_722;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter42_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter43_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter44_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter45_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter46_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter47_reg;
    reg   [63:0] add_i1_1_0_3_reg_722_pp0_iter48_reg;
    wire   [63:0] grp_fu_116_p2;
    reg   [63:0] add_i1_1_1_2_reg_728;
    wire   [63:0] grp_fu_120_p2;
    reg   [63:0] add_i1_1_2_2_reg_733;
    wire   [63:0] grp_fu_124_p2;
    reg   [63:0] add_i1_1_3_2_reg_738;
    wire   [63:0] grp_fu_128_p2;
    reg   [63:0] add_i1_2_0_3_reg_743;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter42_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter43_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter44_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter45_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter46_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter47_reg;
    reg   [63:0] add_i1_2_0_3_reg_743_pp0_iter48_reg;
    wire   [63:0] grp_fu_132_p2;
    reg   [63:0] add_i1_2_1_2_reg_749;
    wire   [63:0] grp_fu_136_p2;
    reg   [63:0] add_i1_2_2_2_reg_754;
    wire   [63:0] grp_fu_140_p2;
    reg   [63:0] add_i1_2_3_2_reg_759;
    wire   [63:0] grp_fu_144_p2;
    reg   [63:0] add_i1_0_1_3_reg_764;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter49_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter50_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter51_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter52_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter53_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter54_reg;
    reg   [63:0] add_i1_0_1_3_reg_764_pp0_iter55_reg;
    wire   [63:0] grp_fu_148_p2;
    reg   [63:0] add_i1_0_2_3_reg_771;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter49_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter50_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter51_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter52_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter53_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter54_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter55_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter56_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter57_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter58_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter59_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter60_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter61_reg;
    reg   [63:0] add_i1_0_2_3_reg_771_pp0_iter62_reg;
    wire   [63:0] grp_fu_152_p2;
    reg   [63:0] add_i1_0_3_3_reg_777;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter49_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter50_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter51_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter52_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter53_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter54_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter55_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter56_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter57_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter58_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter59_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter60_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter61_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter62_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter63_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter64_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter65_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter66_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter67_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter68_reg;
    reg   [63:0] add_i1_0_3_3_reg_777_pp0_iter69_reg;
    wire   [63:0] grp_fu_156_p2;
    reg   [63:0] add_i1_1_1_3_reg_783;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter49_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter50_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter51_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter52_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter53_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter54_reg;
    reg   [63:0] add_i1_1_1_3_reg_783_pp0_iter55_reg;
    wire   [63:0] grp_fu_160_p2;
    reg   [63:0] add_i1_1_2_3_reg_790;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter49_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter50_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter51_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter52_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter53_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter54_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter55_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter56_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter57_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter58_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter59_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter60_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter61_reg;
    reg   [63:0] add_i1_1_2_3_reg_790_pp0_iter62_reg;
    wire   [63:0] grp_fu_164_p2;
    reg   [63:0] add_i1_1_3_3_reg_796;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter49_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter50_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter51_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter52_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter53_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter54_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter55_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter56_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter57_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter58_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter59_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter60_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter61_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter62_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter63_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter64_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter65_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter66_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter67_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter68_reg;
    reg   [63:0] add_i1_1_3_3_reg_796_pp0_iter69_reg;
    wire   [63:0] grp_fu_168_p2;
    reg   [63:0] add_i1_2_1_3_reg_802;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter49_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter50_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter51_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter52_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter53_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter54_reg;
    reg   [63:0] add_i1_2_1_3_reg_802_pp0_iter55_reg;
    wire   [63:0] grp_fu_172_p2;
    reg   [63:0] add_i1_2_2_3_reg_809;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter49_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter50_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter51_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter52_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter53_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter54_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter55_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter56_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter57_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter58_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter59_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter60_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter61_reg;
    reg   [63:0] add_i1_2_2_3_reg_809_pp0_iter62_reg;
    wire   [63:0] grp_fu_176_p2;
    reg   [63:0] add_i1_2_3_3_reg_815;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter49_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter50_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter51_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter52_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter53_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter54_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter55_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter56_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter57_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter58_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter59_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter60_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter61_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter62_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter63_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter64_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter65_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter66_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter67_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter68_reg;
    reg   [63:0] add_i1_2_3_3_reg_815_pp0_iter69_reg;
    wire   [63:0] grp_fu_385_p2;
    reg   [63:0] mul_i2_0_1_reg_821;
    wire   [63:0] grp_fu_390_p2;
    reg   [63:0] mul_i2_1_1_reg_826;
    wire   [63:0] grp_fu_395_p2;
    reg   [63:0] mul_i2_2_1_reg_831;
    wire   [63:0] grp_fu_180_p2;
    reg   [63:0] add_i2_reg_836;
    wire   [63:0] grp_fu_400_p2;
    reg   [63:0] mul_i2_0_0_1_reg_841;
    wire   [63:0] grp_fu_185_p2;
    reg   [63:0] add_i2_0_1_reg_847;
    wire   [63:0] grp_fu_405_p2;
    reg   [63:0] mul_i2_0_2_1_reg_854;
    wire   [63:0] grp_fu_190_p2;
    reg   [63:0] add_i2_1_reg_859;
    wire   [63:0] grp_fu_410_p2;
    reg   [63:0] mul_i2_1_0_1_reg_864;
    wire   [63:0] grp_fu_195_p2;
    reg   [63:0] add_i2_1_1_reg_870;
    wire   [63:0] grp_fu_415_p2;
    reg   [63:0] mul_i2_1_2_1_reg_877;
    wire   [63:0] grp_fu_200_p2;
    reg   [63:0] add_i2_2_reg_882;
    wire   [63:0] grp_fu_420_p2;
    reg   [63:0] mul_i2_2_0_1_reg_887;
    wire   [63:0] grp_fu_205_p2;
    reg   [63:0] add_i2_2_1_reg_893;
    wire   [63:0] grp_fu_425_p2;
    reg   [63:0] mul_i2_2_2_1_reg_900;
    wire   [63:0] grp_fu_210_p2;
    reg   [63:0] add_i2_0_0_1_reg_905;
    wire   [63:0] grp_fu_430_p2;
    reg   [63:0] mul_i2_0_0_2_reg_910;
    wire   [63:0] grp_fu_214_p2;
    reg   [63:0] add_i2_0_1_1_reg_917;
    wire   [63:0] grp_fu_218_p2;
    reg   [63:0] add_i2_0_2_1_reg_922;
    wire   [63:0] grp_fu_222_p2;
    reg   [63:0] add_i2_0_3_1_reg_927;
    wire   [63:0] grp_fu_226_p2;
    reg   [63:0] add_i2_1_0_1_reg_932;
    wire   [63:0] grp_fu_435_p2;
    reg   [63:0] mul_i2_1_0_2_reg_937;
    wire   [63:0] grp_fu_230_p2;
    reg   [63:0] add_i2_1_1_1_reg_944;
    wire   [63:0] grp_fu_234_p2;
    reg   [63:0] add_i2_1_2_1_reg_949;
    wire   [63:0] grp_fu_238_p2;
    reg   [63:0] add_i2_1_3_1_reg_954;
    wire   [63:0] grp_fu_242_p2;
    reg   [63:0] add_i2_2_0_1_reg_959;
    wire   [63:0] grp_fu_440_p2;
    reg   [63:0] mul_i2_2_0_2_reg_964;
    wire   [63:0] grp_fu_246_p2;
    reg   [63:0] add_i2_2_1_1_reg_971;
    wire   [63:0] grp_fu_250_p2;
    reg   [63:0] add_i2_2_2_1_reg_976;
    wire   [63:0] grp_fu_254_p2;
    reg   [63:0] add_i2_2_3_1_reg_981;
    wire   [63:0] grp_fu_258_p2;
    reg   [63:0] add_i2_0_0_2_reg_986;
    wire   [63:0] grp_fu_445_p2;
    reg   [63:0] mul_i2_0_0_3_reg_991;
    wire   [63:0] grp_fu_262_p2;
    reg   [63:0] add_i2_0_1_2_reg_998;
    wire   [63:0] grp_fu_266_p2;
    reg   [63:0] add_i2_0_2_2_reg_1003;
    wire   [63:0] grp_fu_270_p2;
    reg   [63:0] add_i2_0_3_2_reg_1008;
    wire   [63:0] grp_fu_274_p2;
    reg   [63:0] add_i2_1_0_2_reg_1013;
    wire   [63:0] grp_fu_450_p2;
    reg   [63:0] mul_i2_1_0_3_reg_1018;
    wire   [63:0] grp_fu_278_p2;
    reg   [63:0] add_i2_1_1_2_reg_1025;
    wire   [63:0] grp_fu_282_p2;
    reg   [63:0] add_i2_1_2_2_reg_1030;
    wire   [63:0] grp_fu_286_p2;
    reg   [63:0] add_i2_1_3_2_reg_1035;
    wire   [63:0] grp_fu_290_p2;
    reg   [63:0] add_i2_2_0_2_reg_1040;
    wire   [63:0] grp_fu_455_p2;
    reg   [63:0] mul_i2_2_0_3_reg_1045;
    wire   [63:0] grp_fu_294_p2;
    reg   [63:0] add_i2_2_1_2_reg_1052;
    wire   [63:0] grp_fu_298_p2;
    reg   [63:0] add_i2_2_2_2_reg_1057;
    wire   [63:0] grp_fu_302_p2;
    reg   [63:0] add_i2_2_3_2_reg_1062;
    wire    ap_block_pp0_stage0;
    wire   [63:0] grp_fu_306_p2;
    wire   [63:0] grp_fu_310_p2;
    wire   [63:0] grp_fu_314_p2;
    wire   [63:0] grp_fu_318_p2;
    wire   [63:0] grp_fu_322_p2;
    wire   [63:0] grp_fu_326_p2;
    wire   [63:0] grp_fu_330_p2;
    wire   [63:0] grp_fu_334_p2;
    wire   [63:0] grp_fu_338_p2;
    wire   [63:0] grp_fu_342_p2;
    wire   [63:0] grp_fu_346_p2;
    wire   [63:0] grp_fu_350_p2;
    reg   [63:0] x_int_reg;
    wire    ap_ce_reg;

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U1 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_538),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_18_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U2 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_538),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_23_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U3 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_544),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_28_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U4 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x_read_reg_532_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_33_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U5 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_reg_565),
        .din1(mul_i1_0_0_1_reg_570),
        .ce(1'b1),
        .dout(grp_fu_38_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U6 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_0_1_reg_583),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_42_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U7 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_553_pp0_iter20_reg),
        .din1(mul_i1_0_1_reg_583),
        .ce(1'b1),
        .dout(grp_fu_47_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U8 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_0_0_1_reg_570),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_51_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U9 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_553_pp0_iter20_reg),
        .din1(mul_i1_0_0_1_reg_570),
        .ce(1'b1),
        .dout(grp_fu_56_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U10 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_1_reg_600),
        .din1(mul_i1_0_0_2_reg_605),
        .ce(1'b1),
        .dout(grp_fu_60_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U11 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_611),
        .din1(add_i_0_1_3_reg_553_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_64_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U12 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_611),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_68_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U13 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_1_reg_617),
        .din1(mul_i1_0_0_2_reg_605),
        .ce(1'b1),
        .dout(grp_fu_72_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U14 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_622),
        .din1(add_i_0_0_3_reg_544_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_76_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U15 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_622),
        .din1(mul_i1_0_1_reg_583_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_80_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U16 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_1_reg_630),
        .din1(mul_i1_2_0_2_reg_635),
        .ce(1'b1),
        .dout(grp_fu_84_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U17 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_622),
        .din1(add_i_0_1_3_reg_553_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_88_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U18 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_622),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_92_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U19 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_2_reg_640),
        .din1(mul_i1_0_0_3_reg_645),
        .ce(1'b1),
        .dout(grp_fu_96_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U20 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_1_reg_658),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_100_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U21 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_663),
        .din1(add_i_0_1_3_reg_553_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_104_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U22 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_663),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_108_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U23 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_2_reg_669),
        .din1(mul_i1_0_0_3_reg_645),
        .ce(1'b1),
        .dout(grp_fu_112_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U24 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_1_reg_674),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_116_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U25 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_679),
        .din1(add_i_0_1_3_reg_553_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_120_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U26 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_679),
        .din1(mul_i1_0_0_1_reg_570_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_124_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U27 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_2_reg_685),
        .din1(mul_i1_0_0_3_reg_645),
        .ce(1'b1),
        .dout(grp_fu_128_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U28 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_1_reg_690),
        .din1(mul_i1_0_1_reg_583_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_132_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U29 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_695),
        .din1(add_i_0_0_3_reg_544_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_136_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U30 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_695),
        .din1(mul_i1_0_1_reg_583_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_140_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U31 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_2_reg_707),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_144_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U32 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_2_reg_712),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_148_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U33 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_2_reg_717),
        .din1(add_i_0_3_3_reg_592_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_152_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U34 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_2_reg_728),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_156_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U35 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_2_reg_733),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_160_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U36 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_2_reg_738),
        .din1(add_i_0_3_3_reg_592_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_164_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U37 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_2_reg_749),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_168_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U38 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_2_reg_754),
        .din1(mul_i1_0_0_3_reg_645_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_172_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U39 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_2_reg_759),
        .din1(add_i_0_3_3_reg_592_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_176_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U40 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_701_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_180_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U41 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_0_1_reg_821),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_185_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U42 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_722_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_190_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U43 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_1_1_reg_826),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_195_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U44 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_743_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_200_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U45 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_2_1_reg_831),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_205_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U46 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_reg_836),
        .din1(mul_i2_0_0_1_reg_841),
        .ce(1'b1),
        .dout(grp_fu_210_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U47 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_847),
        .din1(add_i1_0_1_3_reg_764_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_214_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U48 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_847),
        .din1(mul_i2_0_2_1_reg_854),
        .ce(1'b1),
        .dout(grp_fu_218_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U49 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_847),
        .din1(mul_i2_0_0_1_reg_841),
        .ce(1'b1),
        .dout(grp_fu_222_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U50 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_reg_859),
        .din1(mul_i2_1_0_1_reg_864),
        .ce(1'b1),
        .dout(grp_fu_226_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U51 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_870),
        .din1(add_i1_1_1_3_reg_783_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_230_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U52 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_870),
        .din1(mul_i2_1_2_1_reg_877),
        .ce(1'b1),
        .dout(grp_fu_234_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U53 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_870),
        .din1(mul_i2_1_0_1_reg_864),
        .ce(1'b1),
        .dout(grp_fu_238_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U54 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_reg_882),
        .din1(mul_i2_2_0_1_reg_887),
        .ce(1'b1),
        .dout(grp_fu_242_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U55 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_893),
        .din1(add_i1_2_1_3_reg_802_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_246_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U56 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_893),
        .din1(mul_i2_2_2_1_reg_900),
        .ce(1'b1),
        .dout(grp_fu_250_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U57 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_893),
        .din1(mul_i2_2_0_1_reg_887),
        .ce(1'b1),
        .dout(grp_fu_254_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U58 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_1_reg_905),
        .din1(mul_i2_0_0_2_reg_910),
        .ce(1'b1),
        .dout(grp_fu_258_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U59 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_1_reg_917),
        .din1(mul_i2_0_0_2_reg_910),
        .ce(1'b1),
        .dout(grp_fu_262_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U60 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_1_reg_922),
        .din1(add_i1_0_2_3_reg_771_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_266_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U61 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_1_reg_927),
        .din1(mul_i2_0_0_2_reg_910),
        .ce(1'b1),
        .dout(grp_fu_270_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U62 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_1_reg_932),
        .din1(mul_i2_1_0_2_reg_937),
        .ce(1'b1),
        .dout(grp_fu_274_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U63 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_1_reg_944),
        .din1(mul_i2_1_0_2_reg_937),
        .ce(1'b1),
        .dout(grp_fu_278_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U64 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_1_reg_949),
        .din1(add_i1_1_2_3_reg_790_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_282_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U65 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_1_reg_954),
        .din1(mul_i2_1_0_2_reg_937),
        .ce(1'b1),
        .dout(grp_fu_286_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U66 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_1_reg_959),
        .din1(mul_i2_2_0_2_reg_964),
        .ce(1'b1),
        .dout(grp_fu_290_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U67 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_1_reg_971),
        .din1(mul_i2_2_0_2_reg_964),
        .ce(1'b1),
        .dout(grp_fu_294_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U68 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_1_reg_976),
        .din1(add_i1_2_2_3_reg_809_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_298_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U69 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_1_reg_981),
        .din1(mul_i2_2_0_2_reg_964),
        .ce(1'b1),
        .dout(grp_fu_302_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U70 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_2_reg_986),
        .din1(mul_i2_0_0_3_reg_991),
        .ce(1'b1),
        .dout(grp_fu_306_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U71 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_2_reg_998),
        .din1(mul_i2_0_0_3_reg_991),
        .ce(1'b1),
        .dout(grp_fu_310_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U72 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_2_reg_1003),
        .din1(mul_i2_0_0_3_reg_991),
        .ce(1'b1),
        .dout(grp_fu_314_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U73 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_2_reg_1008),
        .din1(add_i1_0_3_3_reg_777_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_318_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U74 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_2_reg_1013),
        .din1(mul_i2_1_0_3_reg_1018),
        .ce(1'b1),
        .dout(grp_fu_322_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U75 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_2_reg_1025),
        .din1(mul_i2_1_0_3_reg_1018),
        .ce(1'b1),
        .dout(grp_fu_326_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U76 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_2_reg_1030),
        .din1(mul_i2_1_0_3_reg_1018),
        .ce(1'b1),
        .dout(grp_fu_330_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U77 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_2_reg_1035),
        .din1(add_i1_1_3_3_reg_796_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_334_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U78 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_2_reg_1040),
        .din1(mul_i2_2_0_3_reg_1045),
        .ce(1'b1),
        .dout(grp_fu_338_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U79 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_2_reg_1052),
        .din1(mul_i2_2_0_3_reg_1045),
        .ce(1'b1),
        .dout(grp_fu_342_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U80 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_2_reg_1057),
        .din1(mul_i2_2_0_3_reg_1045),
        .ce(1'b1),
        .dout(grp_fu_346_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U81 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_2_reg_1062),
        .din1(add_i1_2_3_3_reg_815_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_350_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U82 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x_int_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_354_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U83 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_553),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_360_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U84 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_544),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_365_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U85 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_553_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_370_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U86 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_544_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_375_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U87 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_3_3_reg_592),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_380_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U88 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_701),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_385_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U89 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_722),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_390_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U90 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_743),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_395_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U91 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_764),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_400_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U92 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_764),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_405_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U93 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_783),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_410_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U94 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_783),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_415_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U95 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_802),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_420_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U96 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_802),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_425_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U97 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_3_reg_771_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_430_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U98 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_3_reg_790_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_435_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U99 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_3_reg_809_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_440_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U100 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_3_reg_777_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_445_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U101 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_3_reg_796_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_450_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U102 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_3_reg_815_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_455_p2)
    );

    always @(posedge ap_clk) begin
        x_int_reg <= x;
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            add_i1_0_0_1_reg_600 <= grp_fu_38_p2;
            add_i1_0_0_2_reg_640 <= grp_fu_60_p2;
            add_i1_0_0_3_reg_701 <= grp_fu_96_p2;
            add_i1_0_0_3_reg_701_pp0_iter42_reg <= add_i1_0_0_3_reg_701;
            add_i1_0_0_3_reg_701_pp0_iter43_reg <= add_i1_0_0_3_reg_701_pp0_iter42_reg;
            add_i1_0_0_3_reg_701_pp0_iter44_reg <= add_i1_0_0_3_reg_701_pp0_iter43_reg;
            add_i1_0_0_3_reg_701_pp0_iter45_reg <= add_i1_0_0_3_reg_701_pp0_iter44_reg;
            add_i1_0_0_3_reg_701_pp0_iter46_reg <= add_i1_0_0_3_reg_701_pp0_iter45_reg;
            add_i1_0_0_3_reg_701_pp0_iter47_reg <= add_i1_0_0_3_reg_701_pp0_iter46_reg;
            add_i1_0_0_3_reg_701_pp0_iter48_reg <= add_i1_0_0_3_reg_701_pp0_iter47_reg;
            add_i1_0_1_1_reg_658 <= grp_fu_64_p2;
            add_i1_0_1_2_reg_707 <= grp_fu_100_p2;
            add_i1_0_1_3_reg_764 <= grp_fu_144_p2;
            add_i1_0_1_3_reg_764_pp0_iter49_reg <= add_i1_0_1_3_reg_764;
            add_i1_0_1_3_reg_764_pp0_iter50_reg <= add_i1_0_1_3_reg_764_pp0_iter49_reg;
            add_i1_0_1_3_reg_764_pp0_iter51_reg <= add_i1_0_1_3_reg_764_pp0_iter50_reg;
            add_i1_0_1_3_reg_764_pp0_iter52_reg <= add_i1_0_1_3_reg_764_pp0_iter51_reg;
            add_i1_0_1_3_reg_764_pp0_iter53_reg <= add_i1_0_1_3_reg_764_pp0_iter52_reg;
            add_i1_0_1_3_reg_764_pp0_iter54_reg <= add_i1_0_1_3_reg_764_pp0_iter53_reg;
            add_i1_0_1_3_reg_764_pp0_iter55_reg <= add_i1_0_1_3_reg_764_pp0_iter54_reg;
            add_i1_0_1_reg_611 <= grp_fu_42_p2;
            add_i1_0_2_1_reg_663 <= grp_fu_68_p2;
            add_i1_0_2_2_reg_712 <= grp_fu_104_p2;
            add_i1_0_2_3_reg_771 <= grp_fu_148_p2;
            add_i1_0_2_3_reg_771_pp0_iter49_reg <= add_i1_0_2_3_reg_771;
            add_i1_0_2_3_reg_771_pp0_iter50_reg <= add_i1_0_2_3_reg_771_pp0_iter49_reg;
            add_i1_0_2_3_reg_771_pp0_iter51_reg <= add_i1_0_2_3_reg_771_pp0_iter50_reg;
            add_i1_0_2_3_reg_771_pp0_iter52_reg <= add_i1_0_2_3_reg_771_pp0_iter51_reg;
            add_i1_0_2_3_reg_771_pp0_iter53_reg <= add_i1_0_2_3_reg_771_pp0_iter52_reg;
            add_i1_0_2_3_reg_771_pp0_iter54_reg <= add_i1_0_2_3_reg_771_pp0_iter53_reg;
            add_i1_0_2_3_reg_771_pp0_iter55_reg <= add_i1_0_2_3_reg_771_pp0_iter54_reg;
            add_i1_0_2_3_reg_771_pp0_iter56_reg <= add_i1_0_2_3_reg_771_pp0_iter55_reg;
            add_i1_0_2_3_reg_771_pp0_iter57_reg <= add_i1_0_2_3_reg_771_pp0_iter56_reg;
            add_i1_0_2_3_reg_771_pp0_iter58_reg <= add_i1_0_2_3_reg_771_pp0_iter57_reg;
            add_i1_0_2_3_reg_771_pp0_iter59_reg <= add_i1_0_2_3_reg_771_pp0_iter58_reg;
            add_i1_0_2_3_reg_771_pp0_iter60_reg <= add_i1_0_2_3_reg_771_pp0_iter59_reg;
            add_i1_0_2_3_reg_771_pp0_iter61_reg <= add_i1_0_2_3_reg_771_pp0_iter60_reg;
            add_i1_0_2_3_reg_771_pp0_iter62_reg <= add_i1_0_2_3_reg_771_pp0_iter61_reg;
            add_i1_0_3_2_reg_717 <= grp_fu_108_p2;
            add_i1_0_3_3_reg_777 <= grp_fu_152_p2;
            add_i1_0_3_3_reg_777_pp0_iter49_reg <= add_i1_0_3_3_reg_777;
            add_i1_0_3_3_reg_777_pp0_iter50_reg <= add_i1_0_3_3_reg_777_pp0_iter49_reg;
            add_i1_0_3_3_reg_777_pp0_iter51_reg <= add_i1_0_3_3_reg_777_pp0_iter50_reg;
            add_i1_0_3_3_reg_777_pp0_iter52_reg <= add_i1_0_3_3_reg_777_pp0_iter51_reg;
            add_i1_0_3_3_reg_777_pp0_iter53_reg <= add_i1_0_3_3_reg_777_pp0_iter52_reg;
            add_i1_0_3_3_reg_777_pp0_iter54_reg <= add_i1_0_3_3_reg_777_pp0_iter53_reg;
            add_i1_0_3_3_reg_777_pp0_iter55_reg <= add_i1_0_3_3_reg_777_pp0_iter54_reg;
            add_i1_0_3_3_reg_777_pp0_iter56_reg <= add_i1_0_3_3_reg_777_pp0_iter55_reg;
            add_i1_0_3_3_reg_777_pp0_iter57_reg <= add_i1_0_3_3_reg_777_pp0_iter56_reg;
            add_i1_0_3_3_reg_777_pp0_iter58_reg <= add_i1_0_3_3_reg_777_pp0_iter57_reg;
            add_i1_0_3_3_reg_777_pp0_iter59_reg <= add_i1_0_3_3_reg_777_pp0_iter58_reg;
            add_i1_0_3_3_reg_777_pp0_iter60_reg <= add_i1_0_3_3_reg_777_pp0_iter59_reg;
            add_i1_0_3_3_reg_777_pp0_iter61_reg <= add_i1_0_3_3_reg_777_pp0_iter60_reg;
            add_i1_0_3_3_reg_777_pp0_iter62_reg <= add_i1_0_3_3_reg_777_pp0_iter61_reg;
            add_i1_0_3_3_reg_777_pp0_iter63_reg <= add_i1_0_3_3_reg_777_pp0_iter62_reg;
            add_i1_0_3_3_reg_777_pp0_iter64_reg <= add_i1_0_3_3_reg_777_pp0_iter63_reg;
            add_i1_0_3_3_reg_777_pp0_iter65_reg <= add_i1_0_3_3_reg_777_pp0_iter64_reg;
            add_i1_0_3_3_reg_777_pp0_iter66_reg <= add_i1_0_3_3_reg_777_pp0_iter65_reg;
            add_i1_0_3_3_reg_777_pp0_iter67_reg <= add_i1_0_3_3_reg_777_pp0_iter66_reg;
            add_i1_0_3_3_reg_777_pp0_iter68_reg <= add_i1_0_3_3_reg_777_pp0_iter67_reg;
            add_i1_0_3_3_reg_777_pp0_iter69_reg <= add_i1_0_3_3_reg_777_pp0_iter68_reg;
            add_i1_1_0_1_reg_617 <= grp_fu_47_p2;
            add_i1_1_0_2_reg_669 <= grp_fu_72_p2;
            add_i1_1_0_3_reg_722 <= grp_fu_112_p2;
            add_i1_1_0_3_reg_722_pp0_iter42_reg <= add_i1_1_0_3_reg_722;
            add_i1_1_0_3_reg_722_pp0_iter43_reg <= add_i1_1_0_3_reg_722_pp0_iter42_reg;
            add_i1_1_0_3_reg_722_pp0_iter44_reg <= add_i1_1_0_3_reg_722_pp0_iter43_reg;
            add_i1_1_0_3_reg_722_pp0_iter45_reg <= add_i1_1_0_3_reg_722_pp0_iter44_reg;
            add_i1_1_0_3_reg_722_pp0_iter46_reg <= add_i1_1_0_3_reg_722_pp0_iter45_reg;
            add_i1_1_0_3_reg_722_pp0_iter47_reg <= add_i1_1_0_3_reg_722_pp0_iter46_reg;
            add_i1_1_0_3_reg_722_pp0_iter48_reg <= add_i1_1_0_3_reg_722_pp0_iter47_reg;
            add_i1_1_1_1_reg_674 <= grp_fu_76_p2;
            add_i1_1_1_2_reg_728 <= grp_fu_116_p2;
            add_i1_1_1_3_reg_783 <= grp_fu_156_p2;
            add_i1_1_1_3_reg_783_pp0_iter49_reg <= add_i1_1_1_3_reg_783;
            add_i1_1_1_3_reg_783_pp0_iter50_reg <= add_i1_1_1_3_reg_783_pp0_iter49_reg;
            add_i1_1_1_3_reg_783_pp0_iter51_reg <= add_i1_1_1_3_reg_783_pp0_iter50_reg;
            add_i1_1_1_3_reg_783_pp0_iter52_reg <= add_i1_1_1_3_reg_783_pp0_iter51_reg;
            add_i1_1_1_3_reg_783_pp0_iter53_reg <= add_i1_1_1_3_reg_783_pp0_iter52_reg;
            add_i1_1_1_3_reg_783_pp0_iter54_reg <= add_i1_1_1_3_reg_783_pp0_iter53_reg;
            add_i1_1_1_3_reg_783_pp0_iter55_reg <= add_i1_1_1_3_reg_783_pp0_iter54_reg;
            add_i1_1_1_reg_622 <= grp_fu_51_p2;
            add_i1_1_2_1_reg_679 <= grp_fu_80_p2;
            add_i1_1_2_2_reg_733 <= grp_fu_120_p2;
            add_i1_1_2_3_reg_790 <= grp_fu_160_p2;
            add_i1_1_2_3_reg_790_pp0_iter49_reg <= add_i1_1_2_3_reg_790;
            add_i1_1_2_3_reg_790_pp0_iter50_reg <= add_i1_1_2_3_reg_790_pp0_iter49_reg;
            add_i1_1_2_3_reg_790_pp0_iter51_reg <= add_i1_1_2_3_reg_790_pp0_iter50_reg;
            add_i1_1_2_3_reg_790_pp0_iter52_reg <= add_i1_1_2_3_reg_790_pp0_iter51_reg;
            add_i1_1_2_3_reg_790_pp0_iter53_reg <= add_i1_1_2_3_reg_790_pp0_iter52_reg;
            add_i1_1_2_3_reg_790_pp0_iter54_reg <= add_i1_1_2_3_reg_790_pp0_iter53_reg;
            add_i1_1_2_3_reg_790_pp0_iter55_reg <= add_i1_1_2_3_reg_790_pp0_iter54_reg;
            add_i1_1_2_3_reg_790_pp0_iter56_reg <= add_i1_1_2_3_reg_790_pp0_iter55_reg;
            add_i1_1_2_3_reg_790_pp0_iter57_reg <= add_i1_1_2_3_reg_790_pp0_iter56_reg;
            add_i1_1_2_3_reg_790_pp0_iter58_reg <= add_i1_1_2_3_reg_790_pp0_iter57_reg;
            add_i1_1_2_3_reg_790_pp0_iter59_reg <= add_i1_1_2_3_reg_790_pp0_iter58_reg;
            add_i1_1_2_3_reg_790_pp0_iter60_reg <= add_i1_1_2_3_reg_790_pp0_iter59_reg;
            add_i1_1_2_3_reg_790_pp0_iter61_reg <= add_i1_1_2_3_reg_790_pp0_iter60_reg;
            add_i1_1_2_3_reg_790_pp0_iter62_reg <= add_i1_1_2_3_reg_790_pp0_iter61_reg;
            add_i1_1_3_2_reg_738 <= grp_fu_124_p2;
            add_i1_1_3_3_reg_796 <= grp_fu_164_p2;
            add_i1_1_3_3_reg_796_pp0_iter49_reg <= add_i1_1_3_3_reg_796;
            add_i1_1_3_3_reg_796_pp0_iter50_reg <= add_i1_1_3_3_reg_796_pp0_iter49_reg;
            add_i1_1_3_3_reg_796_pp0_iter51_reg <= add_i1_1_3_3_reg_796_pp0_iter50_reg;
            add_i1_1_3_3_reg_796_pp0_iter52_reg <= add_i1_1_3_3_reg_796_pp0_iter51_reg;
            add_i1_1_3_3_reg_796_pp0_iter53_reg <= add_i1_1_3_3_reg_796_pp0_iter52_reg;
            add_i1_1_3_3_reg_796_pp0_iter54_reg <= add_i1_1_3_3_reg_796_pp0_iter53_reg;
            add_i1_1_3_3_reg_796_pp0_iter55_reg <= add_i1_1_3_3_reg_796_pp0_iter54_reg;
            add_i1_1_3_3_reg_796_pp0_iter56_reg <= add_i1_1_3_3_reg_796_pp0_iter55_reg;
            add_i1_1_3_3_reg_796_pp0_iter57_reg <= add_i1_1_3_3_reg_796_pp0_iter56_reg;
            add_i1_1_3_3_reg_796_pp0_iter58_reg <= add_i1_1_3_3_reg_796_pp0_iter57_reg;
            add_i1_1_3_3_reg_796_pp0_iter59_reg <= add_i1_1_3_3_reg_796_pp0_iter58_reg;
            add_i1_1_3_3_reg_796_pp0_iter60_reg <= add_i1_1_3_3_reg_796_pp0_iter59_reg;
            add_i1_1_3_3_reg_796_pp0_iter61_reg <= add_i1_1_3_3_reg_796_pp0_iter60_reg;
            add_i1_1_3_3_reg_796_pp0_iter62_reg <= add_i1_1_3_3_reg_796_pp0_iter61_reg;
            add_i1_1_3_3_reg_796_pp0_iter63_reg <= add_i1_1_3_3_reg_796_pp0_iter62_reg;
            add_i1_1_3_3_reg_796_pp0_iter64_reg <= add_i1_1_3_3_reg_796_pp0_iter63_reg;
            add_i1_1_3_3_reg_796_pp0_iter65_reg <= add_i1_1_3_3_reg_796_pp0_iter64_reg;
            add_i1_1_3_3_reg_796_pp0_iter66_reg <= add_i1_1_3_3_reg_796_pp0_iter65_reg;
            add_i1_1_3_3_reg_796_pp0_iter67_reg <= add_i1_1_3_3_reg_796_pp0_iter66_reg;
            add_i1_1_3_3_reg_796_pp0_iter68_reg <= add_i1_1_3_3_reg_796_pp0_iter67_reg;
            add_i1_1_3_3_reg_796_pp0_iter69_reg <= add_i1_1_3_3_reg_796_pp0_iter68_reg;
            add_i1_2_0_1_reg_630 <= grp_fu_56_p2;
            add_i1_2_0_2_reg_685 <= grp_fu_84_p2;
            add_i1_2_0_3_reg_743 <= grp_fu_128_p2;
            add_i1_2_0_3_reg_743_pp0_iter42_reg <= add_i1_2_0_3_reg_743;
            add_i1_2_0_3_reg_743_pp0_iter43_reg <= add_i1_2_0_3_reg_743_pp0_iter42_reg;
            add_i1_2_0_3_reg_743_pp0_iter44_reg <= add_i1_2_0_3_reg_743_pp0_iter43_reg;
            add_i1_2_0_3_reg_743_pp0_iter45_reg <= add_i1_2_0_3_reg_743_pp0_iter44_reg;
            add_i1_2_0_3_reg_743_pp0_iter46_reg <= add_i1_2_0_3_reg_743_pp0_iter45_reg;
            add_i1_2_0_3_reg_743_pp0_iter47_reg <= add_i1_2_0_3_reg_743_pp0_iter46_reg;
            add_i1_2_0_3_reg_743_pp0_iter48_reg <= add_i1_2_0_3_reg_743_pp0_iter47_reg;
            add_i1_2_1_1_reg_690 <= grp_fu_88_p2;
            add_i1_2_1_2_reg_749 <= grp_fu_132_p2;
            add_i1_2_1_3_reg_802 <= grp_fu_168_p2;
            add_i1_2_1_3_reg_802_pp0_iter49_reg <= add_i1_2_1_3_reg_802;
            add_i1_2_1_3_reg_802_pp0_iter50_reg <= add_i1_2_1_3_reg_802_pp0_iter49_reg;
            add_i1_2_1_3_reg_802_pp0_iter51_reg <= add_i1_2_1_3_reg_802_pp0_iter50_reg;
            add_i1_2_1_3_reg_802_pp0_iter52_reg <= add_i1_2_1_3_reg_802_pp0_iter51_reg;
            add_i1_2_1_3_reg_802_pp0_iter53_reg <= add_i1_2_1_3_reg_802_pp0_iter52_reg;
            add_i1_2_1_3_reg_802_pp0_iter54_reg <= add_i1_2_1_3_reg_802_pp0_iter53_reg;
            add_i1_2_1_3_reg_802_pp0_iter55_reg <= add_i1_2_1_3_reg_802_pp0_iter54_reg;
            add_i1_2_2_1_reg_695 <= grp_fu_92_p2;
            add_i1_2_2_2_reg_754 <= grp_fu_136_p2;
            add_i1_2_2_3_reg_809 <= grp_fu_172_p2;
            add_i1_2_2_3_reg_809_pp0_iter49_reg <= add_i1_2_2_3_reg_809;
            add_i1_2_2_3_reg_809_pp0_iter50_reg <= add_i1_2_2_3_reg_809_pp0_iter49_reg;
            add_i1_2_2_3_reg_809_pp0_iter51_reg <= add_i1_2_2_3_reg_809_pp0_iter50_reg;
            add_i1_2_2_3_reg_809_pp0_iter52_reg <= add_i1_2_2_3_reg_809_pp0_iter51_reg;
            add_i1_2_2_3_reg_809_pp0_iter53_reg <= add_i1_2_2_3_reg_809_pp0_iter52_reg;
            add_i1_2_2_3_reg_809_pp0_iter54_reg <= add_i1_2_2_3_reg_809_pp0_iter53_reg;
            add_i1_2_2_3_reg_809_pp0_iter55_reg <= add_i1_2_2_3_reg_809_pp0_iter54_reg;
            add_i1_2_2_3_reg_809_pp0_iter56_reg <= add_i1_2_2_3_reg_809_pp0_iter55_reg;
            add_i1_2_2_3_reg_809_pp0_iter57_reg <= add_i1_2_2_3_reg_809_pp0_iter56_reg;
            add_i1_2_2_3_reg_809_pp0_iter58_reg <= add_i1_2_2_3_reg_809_pp0_iter57_reg;
            add_i1_2_2_3_reg_809_pp0_iter59_reg <= add_i1_2_2_3_reg_809_pp0_iter58_reg;
            add_i1_2_2_3_reg_809_pp0_iter60_reg <= add_i1_2_2_3_reg_809_pp0_iter59_reg;
            add_i1_2_2_3_reg_809_pp0_iter61_reg <= add_i1_2_2_3_reg_809_pp0_iter60_reg;
            add_i1_2_2_3_reg_809_pp0_iter62_reg <= add_i1_2_2_3_reg_809_pp0_iter61_reg;
            add_i1_2_3_2_reg_759 <= grp_fu_140_p2;
            add_i1_2_3_3_reg_815 <= grp_fu_176_p2;
            add_i1_2_3_3_reg_815_pp0_iter49_reg <= add_i1_2_3_3_reg_815;
            add_i1_2_3_3_reg_815_pp0_iter50_reg <= add_i1_2_3_3_reg_815_pp0_iter49_reg;
            add_i1_2_3_3_reg_815_pp0_iter51_reg <= add_i1_2_3_3_reg_815_pp0_iter50_reg;
            add_i1_2_3_3_reg_815_pp0_iter52_reg <= add_i1_2_3_3_reg_815_pp0_iter51_reg;
            add_i1_2_3_3_reg_815_pp0_iter53_reg <= add_i1_2_3_3_reg_815_pp0_iter52_reg;
            add_i1_2_3_3_reg_815_pp0_iter54_reg <= add_i1_2_3_3_reg_815_pp0_iter53_reg;
            add_i1_2_3_3_reg_815_pp0_iter55_reg <= add_i1_2_3_3_reg_815_pp0_iter54_reg;
            add_i1_2_3_3_reg_815_pp0_iter56_reg <= add_i1_2_3_3_reg_815_pp0_iter55_reg;
            add_i1_2_3_3_reg_815_pp0_iter57_reg <= add_i1_2_3_3_reg_815_pp0_iter56_reg;
            add_i1_2_3_3_reg_815_pp0_iter58_reg <= add_i1_2_3_3_reg_815_pp0_iter57_reg;
            add_i1_2_3_3_reg_815_pp0_iter59_reg <= add_i1_2_3_3_reg_815_pp0_iter58_reg;
            add_i1_2_3_3_reg_815_pp0_iter60_reg <= add_i1_2_3_3_reg_815_pp0_iter59_reg;
            add_i1_2_3_3_reg_815_pp0_iter61_reg <= add_i1_2_3_3_reg_815_pp0_iter60_reg;
            add_i1_2_3_3_reg_815_pp0_iter62_reg <= add_i1_2_3_3_reg_815_pp0_iter61_reg;
            add_i1_2_3_3_reg_815_pp0_iter63_reg <= add_i1_2_3_3_reg_815_pp0_iter62_reg;
            add_i1_2_3_3_reg_815_pp0_iter64_reg <= add_i1_2_3_3_reg_815_pp0_iter63_reg;
            add_i1_2_3_3_reg_815_pp0_iter65_reg <= add_i1_2_3_3_reg_815_pp0_iter64_reg;
            add_i1_2_3_3_reg_815_pp0_iter66_reg <= add_i1_2_3_3_reg_815_pp0_iter65_reg;
            add_i1_2_3_3_reg_815_pp0_iter67_reg <= add_i1_2_3_3_reg_815_pp0_iter66_reg;
            add_i1_2_3_3_reg_815_pp0_iter68_reg <= add_i1_2_3_3_reg_815_pp0_iter67_reg;
            add_i1_2_3_3_reg_815_pp0_iter69_reg <= add_i1_2_3_3_reg_815_pp0_iter68_reg;
            add_i1_reg_565 <= grp_fu_28_p2;
            add_i2_0_0_1_reg_905 <= grp_fu_210_p2;
            add_i2_0_0_2_reg_986 <= grp_fu_258_p2;
            add_i2_0_1_1_reg_917 <= grp_fu_214_p2;
            add_i2_0_1_2_reg_998 <= grp_fu_262_p2;
            add_i2_0_1_reg_847 <= grp_fu_185_p2;
            add_i2_0_2_1_reg_922 <= grp_fu_218_p2;
            add_i2_0_2_2_reg_1003 <= grp_fu_266_p2;
            add_i2_0_3_1_reg_927 <= grp_fu_222_p2;
            add_i2_0_3_2_reg_1008 <= grp_fu_270_p2;
            add_i2_1_0_1_reg_932 <= grp_fu_226_p2;
            add_i2_1_0_2_reg_1013 <= grp_fu_274_p2;
            add_i2_1_1_1_reg_944 <= grp_fu_230_p2;
            add_i2_1_1_2_reg_1025 <= grp_fu_278_p2;
            add_i2_1_1_reg_870 <= grp_fu_195_p2;
            add_i2_1_2_1_reg_949 <= grp_fu_234_p2;
            add_i2_1_2_2_reg_1030 <= grp_fu_282_p2;
            add_i2_1_3_1_reg_954 <= grp_fu_238_p2;
            add_i2_1_3_2_reg_1035 <= grp_fu_286_p2;
            add_i2_1_reg_859 <= grp_fu_190_p2;
            add_i2_2_0_1_reg_959 <= grp_fu_242_p2;
            add_i2_2_0_2_reg_1040 <= grp_fu_290_p2;
            add_i2_2_1_1_reg_971 <= grp_fu_246_p2;
            add_i2_2_1_2_reg_1052 <= grp_fu_294_p2;
            add_i2_2_1_reg_893 <= grp_fu_205_p2;
            add_i2_2_2_1_reg_976 <= grp_fu_250_p2;
            add_i2_2_2_2_reg_1057 <= grp_fu_298_p2;
            add_i2_2_3_1_reg_981 <= grp_fu_254_p2;
            add_i2_2_3_2_reg_1062 <= grp_fu_302_p2;
            add_i2_2_reg_882 <= grp_fu_200_p2;
            add_i2_reg_836 <= grp_fu_180_p2;
            add_i_0_0_3_reg_544 <= grp_fu_18_p2;
            add_i_0_0_3_reg_544_pp0_iter14_reg <= add_i_0_0_3_reg_544;
            add_i_0_0_3_reg_544_pp0_iter15_reg <= add_i_0_0_3_reg_544_pp0_iter14_reg;
            add_i_0_0_3_reg_544_pp0_iter16_reg <= add_i_0_0_3_reg_544_pp0_iter15_reg;
            add_i_0_0_3_reg_544_pp0_iter17_reg <= add_i_0_0_3_reg_544_pp0_iter16_reg;
            add_i_0_0_3_reg_544_pp0_iter18_reg <= add_i_0_0_3_reg_544_pp0_iter17_reg;
            add_i_0_0_3_reg_544_pp0_iter19_reg <= add_i_0_0_3_reg_544_pp0_iter18_reg;
            add_i_0_0_3_reg_544_pp0_iter20_reg <= add_i_0_0_3_reg_544_pp0_iter19_reg;
            add_i_0_0_3_reg_544_pp0_iter21_reg <= add_i_0_0_3_reg_544_pp0_iter20_reg;
            add_i_0_0_3_reg_544_pp0_iter22_reg <= add_i_0_0_3_reg_544_pp0_iter21_reg;
            add_i_0_0_3_reg_544_pp0_iter23_reg <= add_i_0_0_3_reg_544_pp0_iter22_reg;
            add_i_0_0_3_reg_544_pp0_iter24_reg <= add_i_0_0_3_reg_544_pp0_iter23_reg;
            add_i_0_0_3_reg_544_pp0_iter25_reg <= add_i_0_0_3_reg_544_pp0_iter24_reg;
            add_i_0_0_3_reg_544_pp0_iter26_reg <= add_i_0_0_3_reg_544_pp0_iter25_reg;
            add_i_0_0_3_reg_544_pp0_iter27_reg <= add_i_0_0_3_reg_544_pp0_iter26_reg;
            add_i_0_0_3_reg_544_pp0_iter28_reg <= add_i_0_0_3_reg_544_pp0_iter27_reg;
            add_i_0_0_3_reg_544_pp0_iter29_reg <= add_i_0_0_3_reg_544_pp0_iter28_reg;
            add_i_0_0_3_reg_544_pp0_iter30_reg <= add_i_0_0_3_reg_544_pp0_iter29_reg;
            add_i_0_0_3_reg_544_pp0_iter31_reg <= add_i_0_0_3_reg_544_pp0_iter30_reg;
            add_i_0_0_3_reg_544_pp0_iter32_reg <= add_i_0_0_3_reg_544_pp0_iter31_reg;
            add_i_0_0_3_reg_544_pp0_iter33_reg <= add_i_0_0_3_reg_544_pp0_iter32_reg;
            add_i_0_0_3_reg_544_pp0_iter34_reg <= add_i_0_0_3_reg_544_pp0_iter33_reg;
            add_i_0_1_3_reg_553 <= grp_fu_23_p2;
            add_i_0_1_3_reg_553_pp0_iter14_reg <= add_i_0_1_3_reg_553;
            add_i_0_1_3_reg_553_pp0_iter15_reg <= add_i_0_1_3_reg_553_pp0_iter14_reg;
            add_i_0_1_3_reg_553_pp0_iter16_reg <= add_i_0_1_3_reg_553_pp0_iter15_reg;
            add_i_0_1_3_reg_553_pp0_iter17_reg <= add_i_0_1_3_reg_553_pp0_iter16_reg;
            add_i_0_1_3_reg_553_pp0_iter18_reg <= add_i_0_1_3_reg_553_pp0_iter17_reg;
            add_i_0_1_3_reg_553_pp0_iter19_reg <= add_i_0_1_3_reg_553_pp0_iter18_reg;
            add_i_0_1_3_reg_553_pp0_iter20_reg <= add_i_0_1_3_reg_553_pp0_iter19_reg;
            add_i_0_1_3_reg_553_pp0_iter21_reg <= add_i_0_1_3_reg_553_pp0_iter20_reg;
            add_i_0_1_3_reg_553_pp0_iter22_reg <= add_i_0_1_3_reg_553_pp0_iter21_reg;
            add_i_0_1_3_reg_553_pp0_iter23_reg <= add_i_0_1_3_reg_553_pp0_iter22_reg;
            add_i_0_1_3_reg_553_pp0_iter24_reg <= add_i_0_1_3_reg_553_pp0_iter23_reg;
            add_i_0_1_3_reg_553_pp0_iter25_reg <= add_i_0_1_3_reg_553_pp0_iter24_reg;
            add_i_0_1_3_reg_553_pp0_iter26_reg <= add_i_0_1_3_reg_553_pp0_iter25_reg;
            add_i_0_1_3_reg_553_pp0_iter27_reg <= add_i_0_1_3_reg_553_pp0_iter26_reg;
            add_i_0_1_3_reg_553_pp0_iter28_reg <= add_i_0_1_3_reg_553_pp0_iter27_reg;
            add_i_0_1_3_reg_553_pp0_iter29_reg <= add_i_0_1_3_reg_553_pp0_iter28_reg;
            add_i_0_1_3_reg_553_pp0_iter30_reg <= add_i_0_1_3_reg_553_pp0_iter29_reg;
            add_i_0_1_3_reg_553_pp0_iter31_reg <= add_i_0_1_3_reg_553_pp0_iter30_reg;
            add_i_0_1_3_reg_553_pp0_iter32_reg <= add_i_0_1_3_reg_553_pp0_iter31_reg;
            add_i_0_1_3_reg_553_pp0_iter33_reg <= add_i_0_1_3_reg_553_pp0_iter32_reg;
            add_i_0_1_3_reg_553_pp0_iter34_reg <= add_i_0_1_3_reg_553_pp0_iter33_reg;
            add_i_0_3_3_reg_592 <= grp_fu_33_p2;
            add_i_0_3_3_reg_592_pp0_iter28_reg <= add_i_0_3_3_reg_592;
            add_i_0_3_3_reg_592_pp0_iter29_reg <= add_i_0_3_3_reg_592_pp0_iter28_reg;
            add_i_0_3_3_reg_592_pp0_iter30_reg <= add_i_0_3_3_reg_592_pp0_iter29_reg;
            add_i_0_3_3_reg_592_pp0_iter31_reg <= add_i_0_3_3_reg_592_pp0_iter30_reg;
            add_i_0_3_3_reg_592_pp0_iter32_reg <= add_i_0_3_3_reg_592_pp0_iter31_reg;
            add_i_0_3_3_reg_592_pp0_iter33_reg <= add_i_0_3_3_reg_592_pp0_iter32_reg;
            add_i_0_3_3_reg_592_pp0_iter34_reg <= add_i_0_3_3_reg_592_pp0_iter33_reg;
            add_i_0_3_3_reg_592_pp0_iter35_reg <= add_i_0_3_3_reg_592_pp0_iter34_reg;
            add_i_0_3_3_reg_592_pp0_iter36_reg <= add_i_0_3_3_reg_592_pp0_iter35_reg;
            add_i_0_3_3_reg_592_pp0_iter37_reg <= add_i_0_3_3_reg_592_pp0_iter36_reg;
            add_i_0_3_3_reg_592_pp0_iter38_reg <= add_i_0_3_3_reg_592_pp0_iter37_reg;
            add_i_0_3_3_reg_592_pp0_iter39_reg <= add_i_0_3_3_reg_592_pp0_iter38_reg;
            add_i_0_3_3_reg_592_pp0_iter40_reg <= add_i_0_3_3_reg_592_pp0_iter39_reg;
            add_i_0_3_3_reg_592_pp0_iter41_reg <= add_i_0_3_3_reg_592_pp0_iter40_reg;
            mul_i1_0_0_1_reg_570 <= grp_fu_360_p2;
            mul_i1_0_0_1_reg_570_pp0_iter21_reg <= mul_i1_0_0_1_reg_570;
            mul_i1_0_0_1_reg_570_pp0_iter22_reg <= mul_i1_0_0_1_reg_570_pp0_iter21_reg;
            mul_i1_0_0_1_reg_570_pp0_iter23_reg <= mul_i1_0_0_1_reg_570_pp0_iter22_reg;
            mul_i1_0_0_1_reg_570_pp0_iter24_reg <= mul_i1_0_0_1_reg_570_pp0_iter23_reg;
            mul_i1_0_0_1_reg_570_pp0_iter25_reg <= mul_i1_0_0_1_reg_570_pp0_iter24_reg;
            mul_i1_0_0_1_reg_570_pp0_iter26_reg <= mul_i1_0_0_1_reg_570_pp0_iter25_reg;
            mul_i1_0_0_1_reg_570_pp0_iter27_reg <= mul_i1_0_0_1_reg_570_pp0_iter26_reg;
            mul_i1_0_0_1_reg_570_pp0_iter28_reg <= mul_i1_0_0_1_reg_570_pp0_iter27_reg;
            mul_i1_0_0_1_reg_570_pp0_iter29_reg <= mul_i1_0_0_1_reg_570_pp0_iter28_reg;
            mul_i1_0_0_1_reg_570_pp0_iter30_reg <= mul_i1_0_0_1_reg_570_pp0_iter29_reg;
            mul_i1_0_0_1_reg_570_pp0_iter31_reg <= mul_i1_0_0_1_reg_570_pp0_iter30_reg;
            mul_i1_0_0_1_reg_570_pp0_iter32_reg <= mul_i1_0_0_1_reg_570_pp0_iter31_reg;
            mul_i1_0_0_1_reg_570_pp0_iter33_reg <= mul_i1_0_0_1_reg_570_pp0_iter32_reg;
            mul_i1_0_0_1_reg_570_pp0_iter34_reg <= mul_i1_0_0_1_reg_570_pp0_iter33_reg;
            mul_i1_0_0_2_reg_605 <= grp_fu_370_p2;
            mul_i1_0_0_3_reg_645 <= grp_fu_380_p2;
            mul_i1_0_0_3_reg_645_pp0_iter35_reg <= mul_i1_0_0_3_reg_645;
            mul_i1_0_0_3_reg_645_pp0_iter36_reg <= mul_i1_0_0_3_reg_645_pp0_iter35_reg;
            mul_i1_0_0_3_reg_645_pp0_iter37_reg <= mul_i1_0_0_3_reg_645_pp0_iter36_reg;
            mul_i1_0_0_3_reg_645_pp0_iter38_reg <= mul_i1_0_0_3_reg_645_pp0_iter37_reg;
            mul_i1_0_0_3_reg_645_pp0_iter39_reg <= mul_i1_0_0_3_reg_645_pp0_iter38_reg;
            mul_i1_0_0_3_reg_645_pp0_iter40_reg <= mul_i1_0_0_3_reg_645_pp0_iter39_reg;
            mul_i1_0_0_3_reg_645_pp0_iter41_reg <= mul_i1_0_0_3_reg_645_pp0_iter40_reg;
            mul_i1_0_1_reg_583 <= grp_fu_365_p2;
            mul_i1_0_1_reg_583_pp0_iter21_reg <= mul_i1_0_1_reg_583;
            mul_i1_0_1_reg_583_pp0_iter22_reg <= mul_i1_0_1_reg_583_pp0_iter21_reg;
            mul_i1_0_1_reg_583_pp0_iter23_reg <= mul_i1_0_1_reg_583_pp0_iter22_reg;
            mul_i1_0_1_reg_583_pp0_iter24_reg <= mul_i1_0_1_reg_583_pp0_iter23_reg;
            mul_i1_0_1_reg_583_pp0_iter25_reg <= mul_i1_0_1_reg_583_pp0_iter24_reg;
            mul_i1_0_1_reg_583_pp0_iter26_reg <= mul_i1_0_1_reg_583_pp0_iter25_reg;
            mul_i1_0_1_reg_583_pp0_iter27_reg <= mul_i1_0_1_reg_583_pp0_iter26_reg;
            mul_i1_0_1_reg_583_pp0_iter28_reg <= mul_i1_0_1_reg_583_pp0_iter27_reg;
            mul_i1_0_1_reg_583_pp0_iter29_reg <= mul_i1_0_1_reg_583_pp0_iter28_reg;
            mul_i1_0_1_reg_583_pp0_iter30_reg <= mul_i1_0_1_reg_583_pp0_iter29_reg;
            mul_i1_0_1_reg_583_pp0_iter31_reg <= mul_i1_0_1_reg_583_pp0_iter30_reg;
            mul_i1_0_1_reg_583_pp0_iter32_reg <= mul_i1_0_1_reg_583_pp0_iter31_reg;
            mul_i1_0_1_reg_583_pp0_iter33_reg <= mul_i1_0_1_reg_583_pp0_iter32_reg;
            mul_i1_0_1_reg_583_pp0_iter34_reg <= mul_i1_0_1_reg_583_pp0_iter33_reg;
            mul_i1_2_0_2_reg_635 <= grp_fu_375_p2;
            mul_i2_0_0_1_reg_841 <= grp_fu_400_p2;
            mul_i2_0_0_2_reg_910 <= grp_fu_430_p2;
            mul_i2_0_0_3_reg_991 <= grp_fu_445_p2;
            mul_i2_0_1_reg_821 <= grp_fu_385_p2;
            mul_i2_0_2_1_reg_854 <= grp_fu_405_p2;
            mul_i2_1_0_1_reg_864 <= grp_fu_410_p2;
            mul_i2_1_0_2_reg_937 <= grp_fu_435_p2;
            mul_i2_1_0_3_reg_1018 <= grp_fu_450_p2;
            mul_i2_1_1_reg_826 <= grp_fu_390_p2;
            mul_i2_1_2_1_reg_877 <= grp_fu_415_p2;
            mul_i2_2_0_1_reg_887 <= grp_fu_420_p2;
            mul_i2_2_0_2_reg_964 <= grp_fu_440_p2;
            mul_i2_2_0_3_reg_1045 <= grp_fu_455_p2;
            mul_i2_2_1_reg_831 <= grp_fu_395_p2;
            mul_i2_2_2_1_reg_900 <= grp_fu_425_p2;
            mul_i_0_0_3_reg_538 <= grp_fu_354_p2;
            x_read_reg_532 <= x_int_reg;
            x_read_reg_532_pp0_iter10_reg <= x_read_reg_532_pp0_iter9_reg;
            x_read_reg_532_pp0_iter11_reg <= x_read_reg_532_pp0_iter10_reg;
            x_read_reg_532_pp0_iter12_reg <= x_read_reg_532_pp0_iter11_reg;
            x_read_reg_532_pp0_iter13_reg <= x_read_reg_532_pp0_iter12_reg;
            x_read_reg_532_pp0_iter14_reg <= x_read_reg_532_pp0_iter13_reg;
            x_read_reg_532_pp0_iter15_reg <= x_read_reg_532_pp0_iter14_reg;
            x_read_reg_532_pp0_iter16_reg <= x_read_reg_532_pp0_iter15_reg;
            x_read_reg_532_pp0_iter17_reg <= x_read_reg_532_pp0_iter16_reg;
            x_read_reg_532_pp0_iter18_reg <= x_read_reg_532_pp0_iter17_reg;
            x_read_reg_532_pp0_iter19_reg <= x_read_reg_532_pp0_iter18_reg;
            x_read_reg_532_pp0_iter1_reg <= x_read_reg_532;
            x_read_reg_532_pp0_iter20_reg <= x_read_reg_532_pp0_iter19_reg;
            x_read_reg_532_pp0_iter2_reg <= x_read_reg_532_pp0_iter1_reg;
            x_read_reg_532_pp0_iter3_reg <= x_read_reg_532_pp0_iter2_reg;
            x_read_reg_532_pp0_iter4_reg <= x_read_reg_532_pp0_iter3_reg;
            x_read_reg_532_pp0_iter5_reg <= x_read_reg_532_pp0_iter4_reg;
            x_read_reg_532_pp0_iter6_reg <= x_read_reg_532_pp0_iter5_reg;
            x_read_reg_532_pp0_iter7_reg <= x_read_reg_532_pp0_iter6_reg;
            x_read_reg_532_pp0_iter8_reg <= x_read_reg_532_pp0_iter7_reg;
            x_read_reg_532_pp0_iter9_reg <= x_read_reg_532_pp0_iter8_reg;
        end
    end

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_return_0 = grp_fu_306_p2;

    assign ap_return_1 = grp_fu_310_p2;

    assign ap_return_10 = grp_fu_346_p2;

    assign ap_return_11 = grp_fu_350_p2;

    assign ap_return_2 = grp_fu_314_p2;

    assign ap_return_3 = grp_fu_318_p2;

    assign ap_return_4 = grp_fu_322_p2;

    assign ap_return_5 = grp_fu_326_p2;

    assign ap_return_6 = grp_fu_330_p2;

    assign ap_return_7 = grp_fu_334_p2;

    assign ap_return_8 = grp_fu_338_p2;

    assign ap_return_9 = grp_fu_342_p2;

endmodule  //main_rpyxyzToH_double_2
