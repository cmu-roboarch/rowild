/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_detectCollNode_Pipeline_VITIS_LOOP_276_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    this_cPoints_address0,
    this_cPoints_ce0,
    this_cPoints_we0,
    this_cPoints_d0,
    this_cPoints_address1,
    this_cPoints_ce1,
    this_cPoints_we1,
    this_cPoints_d1,
    this_cAxes_address0,
    this_cAxes_ce0,
    this_cAxes_we0,
    this_cAxes_d0,
    this_TCurr_0_0_address0,
    this_TCurr_0_0_ce0,
    this_TCurr_0_0_q0,
    p_read,
    p_read1,
    p_read2,
    p_read3,
    this_TCurr_0_1_address0,
    this_TCurr_0_1_ce0,
    this_TCurr_0_1_q0,
    p_read16,
    p_read17,
    p_read18,
    p_read19,
    this_TCurr_0_2_address0,
    this_TCurr_0_2_ce0,
    this_TCurr_0_2_q0,
    p_read32,
    p_read33,
    p_read34,
    p_read35,
    this_TCurr_0_3_address0,
    this_TCurr_0_3_ce0,
    this_TCurr_0_3_q0,
    p_read48,
    p_read49,
    p_read50,
    p_read51,
    p_read4,
    p_read5,
    p_read6,
    p_read7,
    p_read20,
    p_read21,
    p_read22,
    p_read23,
    p_read36,
    p_read37,
    p_read38,
    p_read39,
    p_read52,
    p_read53,
    p_read54,
    p_read55,
    p_read8,
    p_read9,
    p_read10,
    p_read11,
    p_read24,
    p_read25,
    p_read26,
    p_read27,
    p_read40,
    p_read41,
    p_read42,
    p_read43,
    p_read56,
    p_read57,
    p_read58,
    p_read59,
    p_read12,
    p_read13,
    p_read14,
    p_read15,
    p_read28,
    p_read29,
    p_read30,
    p_read31,
    p_read44,
    p_read45,
    p_read46,
    p_read47,
    p_read60,
    p_read61,
    p_read62,
    p_read63,
    this_TCurr_1_0_address0,
    this_TCurr_1_0_ce0,
    this_TCurr_1_0_q0,
    this_TCurr_1_1_address0,
    this_TCurr_1_1_ce0,
    this_TCurr_1_1_q0,
    this_TCurr_1_2_address0,
    this_TCurr_1_2_ce0,
    this_TCurr_1_2_q0,
    this_TCurr_1_3_address0,
    this_TCurr_1_3_ce0,
    this_TCurr_1_3_q0,
    this_TCurr_2_0_address0,
    this_TCurr_2_0_ce0,
    this_TCurr_2_0_q0,
    this_TCurr_2_1_address0,
    this_TCurr_2_1_ce0,
    this_TCurr_2_1_q0,
    this_TCurr_2_2_address0,
    this_TCurr_2_2_ce0,
    this_TCurr_2_2_q0,
    this_TCurr_2_3_address0,
    this_TCurr_2_3_ce0,
    this_TCurr_2_3_q0,
    l_TColl_0_0_0_constprop_i,
    l_TColl_0_0_0_constprop_o,
    l_TColl_0_0_0_constprop_o_ap_vld,
    l_TColl_0_0_1_constprop_i,
    l_TColl_0_0_1_constprop_o,
    l_TColl_0_0_1_constprop_o_ap_vld,
    l_TColl_0_0_2_constprop_i,
    l_TColl_0_0_2_constprop_o,
    l_TColl_0_0_2_constprop_o_ap_vld,
    l_TColl_0_0_3_constprop_i,
    l_TColl_0_0_3_constprop_o,
    l_TColl_0_0_3_constprop_o_ap_vld,
    l_TColl_1_0_0_constprop_i,
    l_TColl_1_0_0_constprop_o,
    l_TColl_1_0_0_constprop_o_ap_vld,
    l_TColl_1_0_1_constprop_i,
    l_TColl_1_0_1_constprop_o,
    l_TColl_1_0_1_constprop_o_ap_vld,
    l_TColl_1_0_2_constprop_i,
    l_TColl_1_0_2_constprop_o,
    l_TColl_1_0_2_constprop_o_ap_vld,
    l_TColl_1_0_3_constprop_i,
    l_TColl_1_0_3_constprop_o,
    l_TColl_1_0_3_constprop_o_ap_vld,
    l_TColl_2_0_0_constprop_i,
    l_TColl_2_0_0_constprop_o,
    l_TColl_2_0_0_constprop_o_ap_vld,
    l_TColl_2_0_1_constprop_i,
    l_TColl_2_0_1_constprop_o,
    l_TColl_2_0_1_constprop_o_ap_vld,
    l_TColl_2_0_2_constprop_i,
    l_TColl_2_0_2_constprop_o,
    l_TColl_2_0_2_constprop_o_ap_vld,
    l_TColl_2_0_3_constprop_i,
    l_TColl_2_0_3_constprop_o,
    l_TColl_2_0_3_constprop_o_ap_vld,
    l_TColl_0_1_0_constprop_i,
    l_TColl_0_1_0_constprop_o,
    l_TColl_0_1_0_constprop_o_ap_vld,
    l_TColl_0_1_1_constprop_i,
    l_TColl_0_1_1_constprop_o,
    l_TColl_0_1_1_constprop_o_ap_vld,
    l_TColl_0_1_2_constprop_i,
    l_TColl_0_1_2_constprop_o,
    l_TColl_0_1_2_constprop_o_ap_vld,
    l_TColl_0_1_3_constprop_i,
    l_TColl_0_1_3_constprop_o,
    l_TColl_0_1_3_constprop_o_ap_vld,
    l_TColl_1_1_0_constprop_i,
    l_TColl_1_1_0_constprop_o,
    l_TColl_1_1_0_constprop_o_ap_vld,
    l_TColl_1_1_1_constprop_i,
    l_TColl_1_1_1_constprop_o,
    l_TColl_1_1_1_constprop_o_ap_vld,
    l_TColl_1_1_2_constprop_i,
    l_TColl_1_1_2_constprop_o,
    l_TColl_1_1_2_constprop_o_ap_vld,
    l_TColl_1_1_3_constprop_i,
    l_TColl_1_1_3_constprop_o,
    l_TColl_1_1_3_constprop_o_ap_vld,
    l_TColl_2_1_0_constprop_i,
    l_TColl_2_1_0_constprop_o,
    l_TColl_2_1_0_constprop_o_ap_vld,
    l_TColl_2_1_1_constprop_i,
    l_TColl_2_1_1_constprop_o,
    l_TColl_2_1_1_constprop_o_ap_vld,
    l_TColl_2_1_2_constprop_i,
    l_TColl_2_1_2_constprop_o,
    l_TColl_2_1_2_constprop_o_ap_vld,
    l_TColl_2_1_3_constprop_i,
    l_TColl_2_1_3_constprop_o,
    l_TColl_2_1_3_constprop_o_ap_vld,
    l_TColl_0_2_0_constprop_i,
    l_TColl_0_2_0_constprop_o,
    l_TColl_0_2_0_constprop_o_ap_vld,
    l_TColl_0_2_1_constprop_i,
    l_TColl_0_2_1_constprop_o,
    l_TColl_0_2_1_constprop_o_ap_vld,
    l_TColl_0_2_2_constprop_i,
    l_TColl_0_2_2_constprop_o,
    l_TColl_0_2_2_constprop_o_ap_vld,
    l_TColl_0_2_3_constprop_i,
    l_TColl_0_2_3_constprop_o,
    l_TColl_0_2_3_constprop_o_ap_vld,
    l_TColl_1_2_0_constprop_i,
    l_TColl_1_2_0_constprop_o,
    l_TColl_1_2_0_constprop_o_ap_vld,
    l_TColl_1_2_1_constprop_i,
    l_TColl_1_2_1_constprop_o,
    l_TColl_1_2_1_constprop_o_ap_vld,
    l_TColl_1_2_2_constprop_i,
    l_TColl_1_2_2_constprop_o,
    l_TColl_1_2_2_constprop_o_ap_vld,
    l_TColl_1_2_3_constprop_i,
    l_TColl_1_2_3_constprop_o,
    l_TColl_1_2_3_constprop_o_ap_vld,
    l_TColl_2_2_0_constprop_i,
    l_TColl_2_2_0_constprop_o,
    l_TColl_2_2_0_constprop_o_ap_vld,
    l_TColl_2_2_1_constprop_i,
    l_TColl_2_2_1_constprop_o,
    l_TColl_2_2_1_constprop_o_ap_vld,
    l_TColl_2_2_2_constprop_i,
    l_TColl_2_2_2_constprop_o,
    l_TColl_2_2_2_constprop_o_ap_vld,
    l_TColl_2_2_3_constprop_i,
    l_TColl_2_2_3_constprop_o,
    l_TColl_2_2_3_constprop_o_ap_vld,
    l_TColl_0_3_0_constprop_i,
    l_TColl_0_3_0_constprop_o,
    l_TColl_0_3_0_constprop_o_ap_vld,
    l_TColl_0_3_1_constprop_i,
    l_TColl_0_3_1_constprop_o,
    l_TColl_0_3_1_constprop_o_ap_vld,
    l_TColl_0_3_2_constprop_i,
    l_TColl_0_3_2_constprop_o,
    l_TColl_0_3_2_constprop_o_ap_vld,
    l_TColl_0_3_3_constprop_i,
    l_TColl_0_3_3_constprop_o,
    l_TColl_0_3_3_constprop_o_ap_vld,
    l_TColl_1_3_0_constprop_i,
    l_TColl_1_3_0_constprop_o,
    l_TColl_1_3_0_constprop_o_ap_vld,
    l_TColl_1_3_1_constprop_i,
    l_TColl_1_3_1_constprop_o,
    l_TColl_1_3_1_constprop_o_ap_vld,
    l_TColl_1_3_2_constprop_i,
    l_TColl_1_3_2_constprop_o,
    l_TColl_1_3_2_constprop_o_ap_vld,
    l_TColl_1_3_3_constprop_i,
    l_TColl_1_3_3_constprop_o,
    l_TColl_1_3_3_constprop_o_ap_vld,
    l_TColl_2_3_0_constprop_i,
    l_TColl_2_3_0_constprop_o,
    l_TColl_2_3_0_constprop_o_ap_vld,
    l_TColl_2_3_1_constprop_i,
    l_TColl_2_3_1_constprop_o,
    l_TColl_2_3_1_constprop_o_ap_vld,
    l_TColl_2_3_2_constprop_i,
    l_TColl_2_3_2_constprop_o,
    l_TColl_2_3_2_constprop_o_ap_vld,
    l_TColl_2_3_3_constprop_i,
    l_TColl_2_3_3_constprop_o,
    l_TColl_2_3_3_constprop_o_ap_vld,
    grp_fu_1754_p_din0,
    grp_fu_1754_p_din1,
    grp_fu_1754_p_opcode,
    grp_fu_1754_p_dout0,
    grp_fu_1754_p_ce,
    grp_fu_1758_p_din0,
    grp_fu_1758_p_din1,
    grp_fu_1758_p_dout0,
    grp_fu_1758_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 53'd1;
    parameter ap_ST_fsm_pp0_stage1 = 53'd2;
    parameter ap_ST_fsm_pp0_stage2 = 53'd4;
    parameter ap_ST_fsm_pp0_stage3 = 53'd8;
    parameter ap_ST_fsm_pp0_stage4 = 53'd16;
    parameter ap_ST_fsm_pp0_stage5 = 53'd32;
    parameter ap_ST_fsm_pp0_stage6 = 53'd64;
    parameter ap_ST_fsm_pp0_stage7 = 53'd128;
    parameter ap_ST_fsm_pp0_stage8 = 53'd256;
    parameter ap_ST_fsm_pp0_stage9 = 53'd512;
    parameter ap_ST_fsm_pp0_stage10 = 53'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 53'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 53'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 53'd8192;
    parameter ap_ST_fsm_pp0_stage14 = 53'd16384;
    parameter ap_ST_fsm_pp0_stage15 = 53'd32768;
    parameter ap_ST_fsm_pp0_stage16 = 53'd65536;
    parameter ap_ST_fsm_pp0_stage17 = 53'd131072;
    parameter ap_ST_fsm_pp0_stage18 = 53'd262144;
    parameter ap_ST_fsm_pp0_stage19 = 53'd524288;
    parameter ap_ST_fsm_pp0_stage20 = 53'd1048576;
    parameter ap_ST_fsm_pp0_stage21 = 53'd2097152;
    parameter ap_ST_fsm_pp0_stage22 = 53'd4194304;
    parameter ap_ST_fsm_pp0_stage23 = 53'd8388608;
    parameter ap_ST_fsm_pp0_stage24 = 53'd16777216;
    parameter ap_ST_fsm_pp0_stage25 = 53'd33554432;
    parameter ap_ST_fsm_pp0_stage26 = 53'd67108864;
    parameter ap_ST_fsm_pp0_stage27 = 53'd134217728;
    parameter ap_ST_fsm_pp0_stage28 = 53'd268435456;
    parameter ap_ST_fsm_pp0_stage29 = 53'd536870912;
    parameter ap_ST_fsm_pp0_stage30 = 53'd1073741824;
    parameter ap_ST_fsm_pp0_stage31 = 53'd2147483648;
    parameter ap_ST_fsm_pp0_stage32 = 53'd4294967296;
    parameter ap_ST_fsm_pp0_stage33 = 53'd8589934592;
    parameter ap_ST_fsm_pp0_stage34 = 53'd17179869184;
    parameter ap_ST_fsm_pp0_stage35 = 53'd34359738368;
    parameter ap_ST_fsm_pp0_stage36 = 53'd68719476736;
    parameter ap_ST_fsm_pp0_stage37 = 53'd137438953472;
    parameter ap_ST_fsm_pp0_stage38 = 53'd274877906944;
    parameter ap_ST_fsm_pp0_stage39 = 53'd549755813888;
    parameter ap_ST_fsm_pp0_stage40 = 53'd1099511627776;
    parameter ap_ST_fsm_pp0_stage41 = 53'd2199023255552;
    parameter ap_ST_fsm_pp0_stage42 = 53'd4398046511104;
    parameter ap_ST_fsm_pp0_stage43 = 53'd8796093022208;
    parameter ap_ST_fsm_pp0_stage44 = 53'd17592186044416;
    parameter ap_ST_fsm_pp0_stage45 = 53'd35184372088832;
    parameter ap_ST_fsm_pp0_stage46 = 53'd70368744177664;
    parameter ap_ST_fsm_pp0_stage47 = 53'd140737488355328;
    parameter ap_ST_fsm_pp0_stage48 = 53'd281474976710656;
    parameter ap_ST_fsm_pp0_stage49 = 53'd562949953421312;
    parameter ap_ST_fsm_pp0_stage50 = 53'd1125899906842624;
    parameter ap_ST_fsm_pp0_stage51 = 53'd2251799813685248;
    parameter ap_ST_fsm_pp0_stage52 = 53'd4503599627370496;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] this_cPoints_address0;
    output this_cPoints_ce0;
    output this_cPoints_we0;
    output [63:0] this_cPoints_d0;
    output [6:0] this_cPoints_address1;
    output this_cPoints_ce1;
    output this_cPoints_we1;
    output [63:0] this_cPoints_d1;
    output [5:0] this_cAxes_address0;
    output this_cAxes_ce0;
    output this_cAxes_we0;
    output [63:0] this_cAxes_d0;
    output [2:0] this_TCurr_0_0_address0;
    output this_TCurr_0_0_ce0;
    input [63:0] this_TCurr_0_0_q0;
    input [63:0] p_read;
    input [63:0] p_read1;
    input [63:0] p_read2;
    input [63:0] p_read3;
    output [2:0] this_TCurr_0_1_address0;
    output this_TCurr_0_1_ce0;
    input [63:0] this_TCurr_0_1_q0;
    input [63:0] p_read16;
    input [63:0] p_read17;
    input [63:0] p_read18;
    input [63:0] p_read19;
    output [2:0] this_TCurr_0_2_address0;
    output this_TCurr_0_2_ce0;
    input [63:0] this_TCurr_0_2_q0;
    input [63:0] p_read32;
    input [63:0] p_read33;
    input [63:0] p_read34;
    input [63:0] p_read35;
    output [2:0] this_TCurr_0_3_address0;
    output this_TCurr_0_3_ce0;
    input [63:0] this_TCurr_0_3_q0;
    input [63:0] p_read48;
    input [63:0] p_read49;
    input [63:0] p_read50;
    input [63:0] p_read51;
    input [63:0] p_read4;
    input [63:0] p_read5;
    input [63:0] p_read6;
    input [63:0] p_read7;
    input [63:0] p_read20;
    input [63:0] p_read21;
    input [63:0] p_read22;
    input [63:0] p_read23;
    input [63:0] p_read36;
    input [63:0] p_read37;
    input [63:0] p_read38;
    input [63:0] p_read39;
    input [63:0] p_read52;
    input [63:0] p_read53;
    input [63:0] p_read54;
    input [63:0] p_read55;
    input [63:0] p_read8;
    input [63:0] p_read9;
    input [63:0] p_read10;
    input [63:0] p_read11;
    input [63:0] p_read24;
    input [63:0] p_read25;
    input [63:0] p_read26;
    input [63:0] p_read27;
    input [63:0] p_read40;
    input [63:0] p_read41;
    input [63:0] p_read42;
    input [63:0] p_read43;
    input [63:0] p_read56;
    input [63:0] p_read57;
    input [63:0] p_read58;
    input [63:0] p_read59;
    input [63:0] p_read12;
    input [63:0] p_read13;
    input [63:0] p_read14;
    input [63:0] p_read15;
    input [63:0] p_read28;
    input [63:0] p_read29;
    input [63:0] p_read30;
    input [63:0] p_read31;
    input [63:0] p_read44;
    input [63:0] p_read45;
    input [63:0] p_read46;
    input [63:0] p_read47;
    input [63:0] p_read60;
    input [63:0] p_read61;
    input [63:0] p_read62;
    input [63:0] p_read63;
    output [2:0] this_TCurr_1_0_address0;
    output this_TCurr_1_0_ce0;
    input [63:0] this_TCurr_1_0_q0;
    output [2:0] this_TCurr_1_1_address0;
    output this_TCurr_1_1_ce0;
    input [63:0] this_TCurr_1_1_q0;
    output [2:0] this_TCurr_1_2_address0;
    output this_TCurr_1_2_ce0;
    input [63:0] this_TCurr_1_2_q0;
    output [2:0] this_TCurr_1_3_address0;
    output this_TCurr_1_3_ce0;
    input [63:0] this_TCurr_1_3_q0;
    output [2:0] this_TCurr_2_0_address0;
    output this_TCurr_2_0_ce0;
    input [63:0] this_TCurr_2_0_q0;
    output [2:0] this_TCurr_2_1_address0;
    output this_TCurr_2_1_ce0;
    input [63:0] this_TCurr_2_1_q0;
    output [2:0] this_TCurr_2_2_address0;
    output this_TCurr_2_2_ce0;
    input [63:0] this_TCurr_2_2_q0;
    output [2:0] this_TCurr_2_3_address0;
    output this_TCurr_2_3_ce0;
    input [63:0] this_TCurr_2_3_q0;
    input [63:0] l_TColl_0_0_0_constprop_i;
    output [63:0] l_TColl_0_0_0_constprop_o;
    output l_TColl_0_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_1_constprop_i;
    output [63:0] l_TColl_0_0_1_constprop_o;
    output l_TColl_0_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_2_constprop_i;
    output [63:0] l_TColl_0_0_2_constprop_o;
    output l_TColl_0_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_3_constprop_i;
    output [63:0] l_TColl_0_0_3_constprop_o;
    output l_TColl_0_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_0_constprop_i;
    output [63:0] l_TColl_1_0_0_constprop_o;
    output l_TColl_1_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_1_constprop_i;
    output [63:0] l_TColl_1_0_1_constprop_o;
    output l_TColl_1_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_2_constprop_i;
    output [63:0] l_TColl_1_0_2_constprop_o;
    output l_TColl_1_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_3_constprop_i;
    output [63:0] l_TColl_1_0_3_constprop_o;
    output l_TColl_1_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_0_constprop_i;
    output [63:0] l_TColl_2_0_0_constprop_o;
    output l_TColl_2_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_1_constprop_i;
    output [63:0] l_TColl_2_0_1_constprop_o;
    output l_TColl_2_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_2_constprop_i;
    output [63:0] l_TColl_2_0_2_constprop_o;
    output l_TColl_2_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_3_constprop_i;
    output [63:0] l_TColl_2_0_3_constprop_o;
    output l_TColl_2_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_0_constprop_i;
    output [63:0] l_TColl_0_1_0_constprop_o;
    output l_TColl_0_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_1_constprop_i;
    output [63:0] l_TColl_0_1_1_constprop_o;
    output l_TColl_0_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_2_constprop_i;
    output [63:0] l_TColl_0_1_2_constprop_o;
    output l_TColl_0_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_3_constprop_i;
    output [63:0] l_TColl_0_1_3_constprop_o;
    output l_TColl_0_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_0_constprop_i;
    output [63:0] l_TColl_1_1_0_constprop_o;
    output l_TColl_1_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_1_constprop_i;
    output [63:0] l_TColl_1_1_1_constprop_o;
    output l_TColl_1_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_2_constprop_i;
    output [63:0] l_TColl_1_1_2_constprop_o;
    output l_TColl_1_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_3_constprop_i;
    output [63:0] l_TColl_1_1_3_constprop_o;
    output l_TColl_1_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_0_constprop_i;
    output [63:0] l_TColl_2_1_0_constprop_o;
    output l_TColl_2_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_1_constprop_i;
    output [63:0] l_TColl_2_1_1_constprop_o;
    output l_TColl_2_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_2_constprop_i;
    output [63:0] l_TColl_2_1_2_constprop_o;
    output l_TColl_2_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_3_constprop_i;
    output [63:0] l_TColl_2_1_3_constprop_o;
    output l_TColl_2_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_0_constprop_i;
    output [63:0] l_TColl_0_2_0_constprop_o;
    output l_TColl_0_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_1_constprop_i;
    output [63:0] l_TColl_0_2_1_constprop_o;
    output l_TColl_0_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_2_constprop_i;
    output [63:0] l_TColl_0_2_2_constprop_o;
    output l_TColl_0_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_3_constprop_i;
    output [63:0] l_TColl_0_2_3_constprop_o;
    output l_TColl_0_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_0_constprop_i;
    output [63:0] l_TColl_1_2_0_constprop_o;
    output l_TColl_1_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_1_constprop_i;
    output [63:0] l_TColl_1_2_1_constprop_o;
    output l_TColl_1_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_2_constprop_i;
    output [63:0] l_TColl_1_2_2_constprop_o;
    output l_TColl_1_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_3_constprop_i;
    output [63:0] l_TColl_1_2_3_constprop_o;
    output l_TColl_1_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_0_constprop_i;
    output [63:0] l_TColl_2_2_0_constprop_o;
    output l_TColl_2_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_1_constprop_i;
    output [63:0] l_TColl_2_2_1_constprop_o;
    output l_TColl_2_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_2_constprop_i;
    output [63:0] l_TColl_2_2_2_constprop_o;
    output l_TColl_2_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_3_constprop_i;
    output [63:0] l_TColl_2_2_3_constprop_o;
    output l_TColl_2_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_0_constprop_i;
    output [63:0] l_TColl_0_3_0_constprop_o;
    output l_TColl_0_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_1_constprop_i;
    output [63:0] l_TColl_0_3_1_constprop_o;
    output l_TColl_0_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_2_constprop_i;
    output [63:0] l_TColl_0_3_2_constprop_o;
    output l_TColl_0_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_3_constprop_i;
    output [63:0] l_TColl_0_3_3_constprop_o;
    output l_TColl_0_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_0_constprop_i;
    output [63:0] l_TColl_1_3_0_constprop_o;
    output l_TColl_1_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_1_constprop_i;
    output [63:0] l_TColl_1_3_1_constprop_o;
    output l_TColl_1_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_2_constprop_i;
    output [63:0] l_TColl_1_3_2_constprop_o;
    output l_TColl_1_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_3_constprop_i;
    output [63:0] l_TColl_1_3_3_constprop_o;
    output l_TColl_1_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_0_constprop_i;
    output [63:0] l_TColl_2_3_0_constprop_o;
    output l_TColl_2_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_1_constprop_i;
    output [63:0] l_TColl_2_3_1_constprop_o;
    output l_TColl_2_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_2_constprop_i;
    output [63:0] l_TColl_2_3_2_constprop_o;
    output l_TColl_2_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_3_constprop_i;
    output [63:0] l_TColl_2_3_3_constprop_o;
    output l_TColl_2_3_3_constprop_o_ap_vld;
    output [63:0] grp_fu_1754_p_din0;
    output [63:0] grp_fu_1754_p_din1;
    output [0:0] grp_fu_1754_p_opcode;
    input [63:0] grp_fu_1754_p_dout0;
    output grp_fu_1754_p_ce;
    output [63:0] grp_fu_1758_p_din0;
    output [63:0] grp_fu_1758_p_din1;
    input [63:0] grp_fu_1758_p_dout0;
    output grp_fu_1758_p_ce;

    reg ap_idle;
    reg[5:0] this_cAxes_address0;
    reg this_cAxes_ce0;
    reg this_cAxes_we0;
    reg[63:0] this_cAxes_d0;
    reg this_TCurr_0_0_ce0;
    reg this_TCurr_0_1_ce0;
    reg this_TCurr_0_2_ce0;
    reg this_TCurr_0_3_ce0;
    reg this_TCurr_1_0_ce0;
    reg this_TCurr_1_1_ce0;
    reg this_TCurr_1_2_ce0;
    reg this_TCurr_1_3_ce0;
    reg this_TCurr_2_0_ce0;
    reg this_TCurr_2_1_ce0;
    reg this_TCurr_2_2_ce0;
    reg this_TCurr_2_3_ce0;
    reg[63:0] l_TColl_0_0_0_constprop_o;
    reg l_TColl_0_0_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_0_1_constprop_o;
    reg l_TColl_0_0_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_0_2_constprop_o;
    reg l_TColl_0_0_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_0_3_constprop_o;
    reg l_TColl_0_0_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_0_0_constprop_o;
    reg l_TColl_1_0_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_0_1_constprop_o;
    reg l_TColl_1_0_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_0_2_constprop_o;
    reg l_TColl_1_0_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_0_3_constprop_o;
    reg l_TColl_1_0_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_0_0_constprop_o;
    reg l_TColl_2_0_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_0_1_constprop_o;
    reg l_TColl_2_0_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_0_2_constprop_o;
    reg l_TColl_2_0_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_0_3_constprop_o;
    reg l_TColl_2_0_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_1_0_constprop_o;
    reg l_TColl_0_1_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_1_1_constprop_o;
    reg l_TColl_0_1_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_1_2_constprop_o;
    reg l_TColl_0_1_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_1_3_constprop_o;
    reg l_TColl_0_1_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_1_0_constprop_o;
    reg l_TColl_1_1_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_1_1_constprop_o;
    reg l_TColl_1_1_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_1_2_constprop_o;
    reg l_TColl_1_1_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_1_3_constprop_o;
    reg l_TColl_1_1_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_1_0_constprop_o;
    reg l_TColl_2_1_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_1_1_constprop_o;
    reg l_TColl_2_1_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_1_2_constprop_o;
    reg l_TColl_2_1_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_1_3_constprop_o;
    reg l_TColl_2_1_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_2_0_constprop_o;
    reg l_TColl_0_2_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_2_1_constprop_o;
    reg l_TColl_0_2_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_2_2_constprop_o;
    reg l_TColl_0_2_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_2_3_constprop_o;
    reg l_TColl_0_2_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_2_0_constprop_o;
    reg l_TColl_1_2_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_2_1_constprop_o;
    reg l_TColl_1_2_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_2_2_constprop_o;
    reg l_TColl_1_2_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_2_3_constprop_o;
    reg l_TColl_1_2_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_2_0_constprop_o;
    reg l_TColl_2_2_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_2_1_constprop_o;
    reg l_TColl_2_2_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_2_2_constprop_o;
    reg l_TColl_2_2_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_2_3_constprop_o;
    reg l_TColl_2_2_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_3_0_constprop_o;
    reg l_TColl_0_3_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_3_1_constprop_o;
    reg l_TColl_0_3_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_3_2_constprop_o;
    reg l_TColl_0_3_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_0_3_3_constprop_o;
    reg l_TColl_0_3_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_3_0_constprop_o;
    reg l_TColl_1_3_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_3_1_constprop_o;
    reg l_TColl_1_3_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_3_2_constprop_o;
    reg l_TColl_1_3_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_1_3_3_constprop_o;
    reg l_TColl_1_3_3_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_3_0_constprop_o;
    reg l_TColl_2_3_0_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_3_1_constprop_o;
    reg l_TColl_2_3_1_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_3_2_constprop_o;
    reg l_TColl_2_3_2_constprop_o_ap_vld;
    reg[63:0] l_TColl_2_3_3_constprop_o;
    reg l_TColl_2_3_3_constprop_o_ap_vld;

    (* fsm_encoding = "none" *) reg   [52:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage52;
    wire    ap_block_pp0_stage52_subdone;
    reg   [0:0] icmp_ln276_reg_2049;
    reg    ap_condition_exit_pp0_iter0_stage52;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    reg   [63:0] reg_1094;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    wire    ap_CS_fsm_pp0_stage18;
    wire    ap_block_pp0_stage18_11001;
    wire    ap_CS_fsm_pp0_stage25;
    wire    ap_block_pp0_stage25_11001;
    wire    ap_CS_fsm_pp0_stage32;
    wire    ap_block_pp0_stage32_11001;
    wire    ap_CS_fsm_pp0_stage39;
    wire    ap_block_pp0_stage39_11001;
    wire    ap_CS_fsm_pp0_stage46;
    wire    ap_block_pp0_stage46_11001;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] reg_1100;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    wire    ap_CS_fsm_pp0_stage19;
    wire    ap_block_pp0_stage19_11001;
    wire    ap_CS_fsm_pp0_stage26;
    wire    ap_block_pp0_stage26_11001;
    wire    ap_CS_fsm_pp0_stage33;
    wire    ap_block_pp0_stage33_11001;
    wire    ap_CS_fsm_pp0_stage40;
    wire    ap_block_pp0_stage40_11001;
    wire    ap_CS_fsm_pp0_stage47;
    wire    ap_block_pp0_stage47_11001;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    reg   [63:0] reg_1106;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_11001;
    wire    ap_CS_fsm_pp0_stage20;
    wire    ap_block_pp0_stage20_11001;
    wire    ap_CS_fsm_pp0_stage27;
    wire    ap_block_pp0_stage27_11001;
    wire    ap_CS_fsm_pp0_stage34;
    wire    ap_block_pp0_stage34_11001;
    wire    ap_CS_fsm_pp0_stage41;
    wire    ap_block_pp0_stage41_11001;
    wire    ap_CS_fsm_pp0_stage48;
    wire    ap_block_pp0_stage48_11001;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [63:0] reg_1112;
    wire    ap_CS_fsm_pp0_stage14;
    wire    ap_block_pp0_stage14_11001;
    wire    ap_CS_fsm_pp0_stage21;
    wire    ap_block_pp0_stage21_11001;
    wire    ap_CS_fsm_pp0_stage28;
    wire    ap_block_pp0_stage28_11001;
    wire    ap_CS_fsm_pp0_stage35;
    wire    ap_block_pp0_stage35_11001;
    wire    ap_CS_fsm_pp0_stage42;
    wire    ap_block_pp0_stage42_11001;
    wire    ap_CS_fsm_pp0_stage49;
    wire    ap_block_pp0_stage49_11001;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    reg   [63:0] reg_1118;
    wire    ap_CS_fsm_pp0_stage15;
    wire    ap_block_pp0_stage15_11001;
    wire    ap_CS_fsm_pp0_stage22;
    wire    ap_block_pp0_stage22_11001;
    wire    ap_CS_fsm_pp0_stage29;
    wire    ap_block_pp0_stage29_11001;
    wire    ap_CS_fsm_pp0_stage36;
    wire    ap_block_pp0_stage36_11001;
    wire    ap_CS_fsm_pp0_stage43;
    wire    ap_block_pp0_stage43_11001;
    wire    ap_CS_fsm_pp0_stage50;
    wire    ap_block_pp0_stage50_11001;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    reg   [63:0] reg_1124;
    wire    ap_CS_fsm_pp0_stage16;
    wire    ap_block_pp0_stage16_11001;
    wire    ap_CS_fsm_pp0_stage23;
    wire    ap_block_pp0_stage23_11001;
    wire    ap_CS_fsm_pp0_stage30;
    wire    ap_block_pp0_stage30_11001;
    wire    ap_CS_fsm_pp0_stage37;
    wire    ap_block_pp0_stage37_11001;
    wire    ap_CS_fsm_pp0_stage44;
    wire    ap_block_pp0_stage44_11001;
    wire    ap_CS_fsm_pp0_stage51;
    wire    ap_block_pp0_stage51_11001;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    reg   [63:0] reg_1130;
    wire    ap_CS_fsm_pp0_stage17;
    wire    ap_block_pp0_stage17_11001;
    wire    ap_CS_fsm_pp0_stage24;
    wire    ap_block_pp0_stage24_11001;
    wire    ap_CS_fsm_pp0_stage31;
    wire    ap_block_pp0_stage31_11001;
    wire    ap_CS_fsm_pp0_stage38;
    wire    ap_block_pp0_stage38_11001;
    wire    ap_CS_fsm_pp0_stage45;
    wire    ap_block_pp0_stage45_11001;
    wire    ap_block_pp0_stage52_11001;
    reg   [63:0] reg_1136;
    reg   [63:0] reg_1142;
    reg   [63:0] reg_1148;
    reg   [63:0] reg_1154;
    reg   [63:0] reg_1159;
    reg   [63:0] reg_1165;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    reg   [63:0] reg_1171;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    reg   [63:0] reg_1177;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    reg   [63:0] reg_1182;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    reg   [63:0] reg_1188;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    reg   [63:0] reg_1194;
    reg   [63:0] reg_1200;
    reg   [2:0] i_10_reg_2042;
    reg   [2:0] i_10_reg_2042_pp0_iter1_reg;
    wire   [0:0] icmp_ln276_fu_1213_p2;
    reg   [0:0] icmp_ln276_reg_2049_pp0_iter1_reg;
    wire   [1:0] trunc_ln276_fu_1219_p1;
    reg   [1:0] trunc_ln276_reg_2053;
    reg   [1:0] trunc_ln276_reg_2053_pp0_iter1_reg;
    wire   [63:0] dc_fu_1223_p6;
    reg   [63:0] dc_reg_2061;
    wire   [63:0] tmp_s_fu_1237_p6;
    reg   [63:0] tmp_s_reg_2066;
    wire   [63:0] tmp_286_fu_1251_p6;
    reg   [63:0] tmp_286_reg_2071;
    wire   [63:0] tmp_287_fu_1265_p6;
    reg   [63:0] tmp_287_reg_2076;
    wire   [63:0] tmp_288_fu_1279_p6;
    reg   [63:0] tmp_288_reg_2081;
    wire   [63:0] tmp_289_fu_1293_p6;
    reg   [63:0] tmp_289_reg_2086;
    wire   [63:0] tmp_290_fu_1307_p6;
    reg   [63:0] tmp_290_reg_2091;
    wire   [63:0] tmp_291_fu_1321_p6;
    reg   [63:0] tmp_291_reg_2096;
    wire   [63:0] tmp_292_fu_1335_p6;
    reg   [63:0] tmp_292_reg_2101;
    wire   [63:0] tmp_293_fu_1349_p6;
    reg   [63:0] tmp_293_reg_2106;
    wire   [63:0] tmp_294_fu_1363_p6;
    reg   [63:0] tmp_294_reg_2111;
    wire   [63:0] tmp_295_fu_1377_p6;
    reg   [63:0] tmp_295_reg_2116;
    wire   [63:0] tmp_296_fu_1391_p6;
    reg   [63:0] tmp_296_reg_2121;
    wire   [63:0] tmp_297_fu_1405_p6;
    reg   [63:0] tmp_297_reg_2126;
    wire   [63:0] tmp_298_fu_1419_p6;
    reg   [63:0] tmp_298_reg_2131;
    wire   [63:0] tmp_299_fu_1433_p6;
    reg   [63:0] tmp_299_reg_2136;
    wire   [63:0] tmp_300_fu_1447_p6;
    reg   [63:0] tmp_300_reg_2141;
    reg   [0:0] xs_sign_reg_2146;
    wire   [136:0] zext_ln15_fu_1496_p1;
    reg   [136:0] zext_ln15_reg_2151;
    wire   [0:0] tmp_25_fu_1510_p3;
    reg   [0:0] tmp_25_reg_2156;
    wire   [136:0] zext_ln18_fu_1540_p1;
    reg   [136:0] zext_ln18_reg_2161;
    reg   [2:0] tmp_45_reg_2166;
    wire   [2:0] val_fu_1574_p3;
    reg   [2:0] val_reg_2171;
    reg   [63:0] this_TCurr_0_0_load_reg_2237;
    reg   [63:0] this_TCurr_0_1_load_reg_2242;
    reg   [63:0] this_TCurr_0_2_load_reg_2247;
    reg   [63:0] this_TCurr_0_3_load_reg_2252;
    reg   [63:0] this_TCurr_1_0_load_reg_2257;
    reg   [63:0] this_TCurr_1_1_load_reg_2262;
    reg   [63:0] this_TCurr_1_2_load_reg_2267;
    reg   [63:0] this_TCurr_1_3_load_reg_2272;
    reg   [63:0] this_TCurr_2_0_load_reg_2277;
    reg   [63:0] this_TCurr_2_1_load_reg_2282;
    reg   [63:0] this_TCurr_2_2_load_reg_2287;
    reg   [63:0] this_TCurr_2_3_load_reg_2292;
    wire   [5:0] tmp_fu_1617_p3;
    reg   [5:0] tmp_reg_2297;
    wire   [63:0] tmp_301_fu_1996_p6;
    reg   [63:0] tmp_301_reg_2309;
    wire   [63:0] tmp_302_fu_2009_p6;
    reg   [63:0] tmp_302_reg_2314;
    wire   [63:0] tmp_303_fu_2022_p6;
    reg   [63:0] tmp_303_reg_2319;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage11_subdone;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_ap_start;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_ap_done;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_ap_idle;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_ap_ready;
    wire   [6:0] grp_blockDescToBoundingBox_double_s_fu_979_corners_address0;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_corners_ce0;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_corners_we0;
    wire   [63:0] grp_blockDescToBoundingBox_double_s_fu_979_corners_d0;
    wire   [6:0] grp_blockDescToBoundingBox_double_s_fu_979_corners_address1;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_corners_ce1;
    wire    grp_blockDescToBoundingBox_double_s_fu_979_corners_we1;
    wire   [63:0] grp_blockDescToBoundingBox_double_s_fu_979_corners_d1;
    reg    grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg;
    wire    ap_block_pp0_stage13;
    wire    ap_block_pp0_stage14;
    wire    ap_block_pp0_stage51;
    wire    ap_block_pp0_stage52;
    wire    ap_block_pp0_stage0;
    wire    ap_block_pp0_stage1;
    wire    ap_block_pp0_stage2;
    wire    ap_block_pp0_stage4;
    wire    ap_block_pp0_stage5;
    wire    ap_block_pp0_stage6;
    wire    ap_block_pp0_stage7;
    wire    ap_block_pp0_stage8;
    wire    ap_block_pp0_stage9;
    wire    ap_block_pp0_stage10;
    wire    ap_block_pp0_stage11;
    wire    ap_block_pp0_stage15;
    wire    ap_block_pp0_stage16;
    wire    ap_block_pp0_stage17;
    wire   [63:0] zext_ln278_fu_1591_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln282_fu_1623_p1;
    wire   [63:0] zext_ln282_3_fu_1633_p1;
    wire   [63:0] zext_ln282_6_fu_1643_p1;
    wire   [63:0] zext_ln282_1_fu_1653_p1;
    wire   [63:0] zext_ln282_4_fu_1663_p1;
    wire   [63:0] zext_ln282_7_fu_1673_p1;
    wire   [63:0] zext_ln282_2_fu_1683_p1;
    wire   [63:0] zext_ln282_5_fu_1693_p1;
    wire   [63:0] zext_ln282_8_fu_1703_p1;
    wire    ap_block_pp0_stage12;
    reg   [2:0] i_fu_358;
    wire   [2:0] add_ln276_fu_1607_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_i_10;
    reg   [63:0] grp_fu_1085_p0;
    reg   [63:0] grp_fu_1085_p1;
    wire    ap_block_pp0_stage18;
    wire    ap_block_pp0_stage19;
    wire    ap_block_pp0_stage20;
    wire    ap_block_pp0_stage21;
    wire    ap_block_pp0_stage22;
    wire    ap_block_pp0_stage23;
    wire    ap_block_pp0_stage24;
    wire    ap_block_pp0_stage25;
    wire    ap_block_pp0_stage26;
    wire    ap_block_pp0_stage27;
    wire    ap_block_pp0_stage28;
    wire    ap_block_pp0_stage29;
    wire    ap_block_pp0_stage30;
    wire    ap_block_pp0_stage31;
    wire    ap_block_pp0_stage32;
    wire    ap_block_pp0_stage33;
    wire    ap_block_pp0_stage34;
    wire    ap_block_pp0_stage35;
    wire    ap_block_pp0_stage36;
    wire    ap_block_pp0_stage37;
    wire    ap_block_pp0_stage38;
    wire    ap_block_pp0_stage39;
    wire    ap_block_pp0_stage40;
    wire    ap_block_pp0_stage41;
    wire    ap_block_pp0_stage42;
    wire    ap_block_pp0_stage43;
    wire    ap_block_pp0_stage44;
    wire    ap_block_pp0_stage45;
    wire    ap_block_pp0_stage46;
    wire    ap_block_pp0_stage47;
    wire    ap_block_pp0_stage48;
    wire    ap_block_pp0_stage49;
    wire    ap_block_pp0_stage50;
    reg   [63:0] grp_fu_1090_p0;
    reg   [63:0] grp_fu_1090_p1;
    wire   [63:0] data_fu_1461_p1;
    wire   [51:0] trunc_ln505_fu_1482_p1;
    wire   [53:0] mantissa_fu_1486_p4;
    wire   [10:0] xs_exp_fu_1472_p4;
    wire   [11:0] zext_ln486_fu_1500_p1;
    wire   [11:0] add_ln486_fu_1504_p2;
    wire   [10:0] sub_ln18_fu_1518_p2;
    wire  signed [11:0] sext_ln18_fu_1524_p1;
    wire   [11:0] select_ln18_fu_1528_p3;
    wire  signed [31:0] sext_ln18_1_fu_1536_p1;
    wire   [136:0] lshr_ln18_fu_1544_p2;
    wire   [136:0] shl_ln18_fu_1560_p2;
    wire   [2:0] tmp_46_fu_1564_p4;
    wire   [2:0] result_2_fu_1580_p2;
    wire   [2:0] result_fu_1585_p3;
    wire   [5:0] add_ln282_2_fu_1628_p2;
    wire   [5:0] add_ln282_5_fu_1638_p2;
    wire   [5:0] add_ln282_fu_1648_p2;
    wire   [5:0] add_ln282_3_fu_1658_p2;
    wire   [5:0] add_ln282_6_fu_1668_p2;
    wire   [5:0] add_ln282_1_fu_1678_p2;
    wire   [5:0] add_ln282_4_fu_1688_p2;
    wire   [5:0] add_ln282_7_fu_1698_p2;
    wire    ap_block_pp0_stage12_00001;
    wire    ap_block_pp0_stage13_00001;
    wire    ap_block_pp0_stage14_00001;
    wire    ap_block_pp0_stage15_00001;
    wire    ap_block_pp0_stage16_00001;
    wire    ap_block_pp0_stage17_00001;
    wire    ap_block_pp0_stage18_00001;
    wire    ap_block_pp0_stage19_00001;
    wire    ap_block_pp0_stage20_00001;
    wire    ap_block_pp0_stage21_00001;
    wire    ap_block_pp0_stage22_00001;
    wire    ap_block_pp0_stage23_00001;
    wire    ap_block_pp0_stage24_00001;
    wire    ap_block_pp0_stage25_00001;
    wire    ap_block_pp0_stage26_00001;
    wire    ap_block_pp0_stage27_00001;
    wire    ap_block_pp0_stage28_00001;
    wire    ap_block_pp0_stage29_00001;
    wire    ap_block_pp0_stage30_00001;
    wire    ap_block_pp0_stage31_00001;
    wire    ap_block_pp0_stage32_00001;
    wire    ap_block_pp0_stage33_00001;
    wire    ap_block_pp0_stage34_00001;
    wire    ap_block_pp0_stage35_00001;
    wire    ap_block_pp0_stage36_00001;
    wire    ap_block_pp0_stage37_00001;
    wire    ap_block_pp0_stage38_00001;
    wire    ap_block_pp0_stage39_00001;
    wire    ap_block_pp0_stage40_00001;
    wire    ap_block_pp0_stage41_00001;
    wire    ap_block_pp0_stage42_00001;
    wire    ap_block_pp0_stage43_00001;
    wire    ap_block_pp0_stage44_00001;
    wire    ap_block_pp0_stage45_00001;
    wire    ap_block_pp0_stage46_00001;
    wire    ap_block_pp0_stage47_00001;
    wire    ap_block_pp0_stage48_00001;
    wire    ap_block_pp0_stage49_00001;
    wire    ap_block_pp0_stage50_00001;
    wire    ap_block_pp0_stage51_00001;
    wire    ap_block_pp0_stage52_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage5_00001;
    wire    ap_block_pp0_stage6_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_condition_exit_pp0_iter1_stage11;
    reg    ap_idle_pp0_0to0;
    reg   [52:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to2;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_block_pp0_stage13_subdone;
    wire    ap_block_pp0_stage14_subdone;
    wire    ap_block_pp0_stage15_subdone;
    wire    ap_block_pp0_stage16_subdone;
    wire    ap_block_pp0_stage17_subdone;
    wire    ap_block_pp0_stage18_subdone;
    wire    ap_block_pp0_stage19_subdone;
    wire    ap_block_pp0_stage20_subdone;
    wire    ap_block_pp0_stage21_subdone;
    wire    ap_block_pp0_stage22_subdone;
    wire    ap_block_pp0_stage23_subdone;
    wire    ap_block_pp0_stage24_subdone;
    wire    ap_block_pp0_stage25_subdone;
    wire    ap_block_pp0_stage26_subdone;
    wire    ap_block_pp0_stage27_subdone;
    wire    ap_block_pp0_stage28_subdone;
    wire    ap_block_pp0_stage29_subdone;
    wire    ap_block_pp0_stage30_subdone;
    wire    ap_block_pp0_stage31_subdone;
    wire    ap_block_pp0_stage32_subdone;
    wire    ap_block_pp0_stage33_subdone;
    wire    ap_block_pp0_stage34_subdone;
    wire    ap_block_pp0_stage35_subdone;
    wire    ap_block_pp0_stage36_subdone;
    wire    ap_block_pp0_stage37_subdone;
    wire    ap_block_pp0_stage38_subdone;
    wire    ap_block_pp0_stage39_subdone;
    wire    ap_block_pp0_stage40_subdone;
    wire    ap_block_pp0_stage41_subdone;
    wire    ap_block_pp0_stage42_subdone;
    wire    ap_block_pp0_stage43_subdone;
    wire    ap_block_pp0_stage44_subdone;
    wire    ap_block_pp0_stage45_subdone;
    wire    ap_block_pp0_stage46_subdone;
    wire    ap_block_pp0_stage47_subdone;
    wire    ap_block_pp0_stage48_subdone;
    wire    ap_block_pp0_stage49_subdone;
    wire    ap_block_pp0_stage50_subdone;
    wire    ap_block_pp0_stage51_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 53'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg = 1'b0;
        #0 i_fu_358 = 3'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_blockDescToBoundingBox_double_s grp_blockDescToBoundingBox_double_s_fu_979 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_blockDescToBoundingBox_double_s_fu_979_ap_start),
        .ap_done(grp_blockDescToBoundingBox_double_s_fu_979_ap_done),
        .ap_idle(grp_blockDescToBoundingBox_double_s_fu_979_ap_idle),
        .ap_ready(grp_blockDescToBoundingBox_double_s_fu_979_ap_ready),
        .H_offset(trunc_ln276_reg_2053_pp0_iter1_reg),
        .dim_0_0_val(tmp_301_reg_2309),
        .dim_0_1_val(tmp_302_reg_2314),
        .dim_0_2_val(tmp_303_reg_2319),
        .corners_address0(grp_blockDescToBoundingBox_double_s_fu_979_corners_address0),
        .corners_ce0(grp_blockDescToBoundingBox_double_s_fu_979_corners_ce0),
        .corners_we0(grp_blockDescToBoundingBox_double_s_fu_979_corners_we0),
        .corners_d0(grp_blockDescToBoundingBox_double_s_fu_979_corners_d0),
        .corners_address1(grp_blockDescToBoundingBox_double_s_fu_979_corners_address1),
        .corners_ce1(grp_blockDescToBoundingBox_double_s_fu_979_corners_ce1),
        .corners_we1(grp_blockDescToBoundingBox_double_s_fu_979_corners_we1),
        .corners_d1(grp_blockDescToBoundingBox_double_s_fu_979_corners_d1),
        .l_TColl_0_0_0_constprop(l_TColl_0_0_0_constprop_i),
        .l_TColl_0_0_1_constprop(l_TColl_0_0_1_constprop_i),
        .l_TColl_0_0_2_constprop(l_TColl_0_0_2_constprop_i),
        .l_TColl_0_0_3_constprop(l_TColl_0_0_3_constprop_i),
        .l_TColl_1_0_0_constprop(l_TColl_1_0_0_constprop_i),
        .l_TColl_1_0_1_constprop(l_TColl_1_0_1_constprop_i),
        .l_TColl_1_0_2_constprop(l_TColl_1_0_2_constprop_i),
        .l_TColl_1_0_3_constprop(l_TColl_1_0_3_constprop_i),
        .l_TColl_2_0_0_constprop(l_TColl_2_0_0_constprop_i),
        .l_TColl_2_0_1_constprop(l_TColl_2_0_1_constprop_i),
        .l_TColl_2_0_2_constprop(l_TColl_2_0_2_constprop_i),
        .l_TColl_2_0_3_constprop(l_TColl_2_0_3_constprop_i),
        .l_TColl_0_1_0_constprop(l_TColl_0_1_0_constprop_i),
        .l_TColl_0_1_1_constprop(l_TColl_0_1_1_constprop_i),
        .l_TColl_0_1_2_constprop(l_TColl_0_1_2_constprop_i),
        .l_TColl_0_1_3_constprop(l_TColl_0_1_3_constprop_i),
        .l_TColl_1_1_0_constprop(l_TColl_1_1_0_constprop_i),
        .l_TColl_1_1_1_constprop(l_TColl_1_1_1_constprop_i),
        .l_TColl_1_1_2_constprop(l_TColl_1_1_2_constprop_i),
        .l_TColl_1_1_3_constprop(l_TColl_1_1_3_constprop_i),
        .l_TColl_2_1_0_constprop(l_TColl_2_1_0_constprop_i),
        .l_TColl_2_1_1_constprop(l_TColl_2_1_1_constprop_i),
        .l_TColl_2_1_2_constprop(l_TColl_2_1_2_constprop_i),
        .l_TColl_2_1_3_constprop(l_TColl_2_1_3_constprop_i),
        .l_TColl_0_2_0_constprop(l_TColl_0_2_0_constprop_i),
        .l_TColl_0_2_1_constprop(l_TColl_0_2_1_constprop_i),
        .l_TColl_0_2_2_constprop(l_TColl_0_2_2_constprop_i),
        .l_TColl_0_2_3_constprop(l_TColl_0_2_3_constprop_i),
        .l_TColl_1_2_0_constprop(l_TColl_1_2_0_constprop_i),
        .l_TColl_1_2_1_constprop(l_TColl_1_2_1_constprop_i),
        .l_TColl_1_2_2_constprop(l_TColl_1_2_2_constprop_i),
        .l_TColl_1_2_3_constprop(l_TColl_1_2_3_constprop_i),
        .l_TColl_2_2_0_constprop(l_TColl_2_2_0_constprop_i),
        .l_TColl_2_2_1_constprop(l_TColl_2_2_1_constprop_i),
        .l_TColl_2_2_2_constprop(l_TColl_2_2_2_constprop_i),
        .l_TColl_2_2_3_constprop(l_TColl_2_2_3_constprop_i),
        .l_TColl_0_3_0_constprop(l_TColl_0_3_0_constprop_i),
        .l_TColl_0_3_1_constprop(l_TColl_0_3_1_constprop_i),
        .l_TColl_0_3_2_constprop(l_TColl_0_3_2_constprop_i),
        .l_TColl_0_3_3_constprop(l_TColl_0_3_3_constprop_i),
        .l_TColl_1_3_0_constprop(l_TColl_1_3_0_constprop_i),
        .l_TColl_1_3_1_constprop(l_TColl_1_3_1_constprop_i),
        .l_TColl_1_3_2_constprop(l_TColl_1_3_2_constprop_i),
        .l_TColl_1_3_3_constprop(l_TColl_1_3_3_constprop_i),
        .l_TColl_2_3_0_constprop(l_TColl_2_3_0_constprop_i),
        .l_TColl_2_3_1_constprop(l_TColl_2_3_1_constprop_i),
        .l_TColl_2_3_2_constprop(l_TColl_2_3_2_constprop_i),
        .l_TColl_2_3_3_constprop(l_TColl_2_3_3_constprop_i)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U948 (
        .din0(64'd4607182418800017408),
        .din1(64'd4611686018427387904),
        .din2(64'd4613937818241073152),
        .din3(64'd4616189618054758400),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(dc_fu_1223_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U949 (
        .din0(p_read),
        .din1(p_read1),
        .din2(p_read2),
        .din3(p_read3),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_s_fu_1237_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U950 (
        .din0(p_read16),
        .din1(p_read17),
        .din2(p_read18),
        .din3(p_read19),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_286_fu_1251_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U951 (
        .din0(p_read32),
        .din1(p_read33),
        .din2(p_read34),
        .din3(p_read35),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_287_fu_1265_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U952 (
        .din0(p_read48),
        .din1(p_read49),
        .din2(p_read50),
        .din3(p_read51),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_288_fu_1279_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U953 (
        .din0(p_read4),
        .din1(p_read5),
        .din2(p_read6),
        .din3(p_read7),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_289_fu_1293_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U954 (
        .din0(p_read20),
        .din1(p_read21),
        .din2(p_read22),
        .din3(p_read23),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_290_fu_1307_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U955 (
        .din0(p_read36),
        .din1(p_read37),
        .din2(p_read38),
        .din3(p_read39),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_291_fu_1321_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U956 (
        .din0(p_read52),
        .din1(p_read53),
        .din2(p_read54),
        .din3(p_read55),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_292_fu_1335_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U957 (
        .din0(p_read8),
        .din1(p_read9),
        .din2(p_read10),
        .din3(p_read11),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_293_fu_1349_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U958 (
        .din0(p_read24),
        .din1(p_read25),
        .din2(p_read26),
        .din3(p_read27),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_294_fu_1363_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U959 (
        .din0(p_read40),
        .din1(p_read41),
        .din2(p_read42),
        .din3(p_read43),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_295_fu_1377_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U960 (
        .din0(p_read56),
        .din1(p_read57),
        .din2(p_read58),
        .din3(p_read59),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_296_fu_1391_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U961 (
        .din0(p_read12),
        .din1(p_read13),
        .din2(p_read14),
        .din3(p_read15),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_297_fu_1405_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U962 (
        .din0(p_read28),
        .din1(p_read29),
        .din2(p_read30),
        .din3(p_read31),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_298_fu_1419_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U963 (
        .din0(p_read44),
        .din1(p_read45),
        .din2(p_read46),
        .din3(p_read47),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_299_fu_1433_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U964 (
        .din0(p_read60),
        .din1(p_read61),
        .din2(p_read62),
        .din3(p_read63),
        .din4(trunc_ln276_fu_1219_p1),
        .dout(tmp_300_fu_1447_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U965 (
        .din0(64'd4587366580439587226),
        .din1(64'd4598175219545276416),
        .din2(64'd4589708452245819884),
        .din3(64'd4592590756007337001),
        .din4(trunc_ln276_reg_2053_pp0_iter1_reg),
        .dout(tmp_301_fu_1996_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U966 (
        .din0(64'd4587366580439587226),
        .din1(64'd4587366580439587226),
        .din2(64'd4590140797810047451),
        .din3(64'd4592590756007337001),
        .din4(trunc_ln276_reg_2053_pp0_iter1_reg),
        .dout(tmp_302_fu_2009_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U967 (
        .din0(64'd4598175219545276416),
        .din1(64'd4587366580439587226),
        .din2(64'd4587366580439587226),
        .din3(64'd4589708452245819884),
        .din4(trunc_ln276_reg_2053_pp0_iter1_reg),
        .dout(tmp_303_fu_2022_p6)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage52),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage11_subdone) & (ap_loop_exit_ready_pp0_iter1_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage52)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage52_subdone) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage11_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                ap_enable_reg_pp0_iter2 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage52_subdone) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg <= 1'b1;
            end else if ((grp_blockDescToBoundingBox_double_s_fu_979_ap_ready == 1'b1)) begin
                grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to0 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter1_stage11))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage52_11001) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            i_fu_358 <= 3'd0;
        end else if (((icmp_ln276_reg_2049 == 1'd0) & (1'b0 == ap_block_pp0_stage52_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
            i_fu_358 <= add_ln276_fu_1607_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            dc_reg_2061 <= dc_fu_1223_p6;
            i_10_reg_2042 <= ap_sig_allocacmp_i_10;
            i_10_reg_2042_pp0_iter1_reg <= i_10_reg_2042;
            icmp_ln276_reg_2049 <= icmp_ln276_fu_1213_p2;
            icmp_ln276_reg_2049_pp0_iter1_reg <= icmp_ln276_reg_2049;
            tmp_286_reg_2071 <= tmp_286_fu_1251_p6;
            tmp_287_reg_2076 <= tmp_287_fu_1265_p6;
            tmp_288_reg_2081 <= tmp_288_fu_1279_p6;
            tmp_289_reg_2086 <= tmp_289_fu_1293_p6;
            tmp_290_reg_2091 <= tmp_290_fu_1307_p6;
            tmp_291_reg_2096 <= tmp_291_fu_1321_p6;
            tmp_292_reg_2101 <= tmp_292_fu_1335_p6;
            tmp_293_reg_2106 <= tmp_293_fu_1349_p6;
            tmp_294_reg_2111 <= tmp_294_fu_1363_p6;
            tmp_295_reg_2116 <= tmp_295_fu_1377_p6;
            tmp_296_reg_2121 <= tmp_296_fu_1391_p6;
            tmp_297_reg_2126 <= tmp_297_fu_1405_p6;
            tmp_298_reg_2131 <= tmp_298_fu_1419_p6;
            tmp_299_reg_2136 <= tmp_299_fu_1433_p6;
            tmp_300_reg_2141 <= tmp_300_fu_1447_p6;
            tmp_s_reg_2066 <= tmp_s_fu_1237_p6;
            trunc_ln276_reg_2053 <= trunc_ln276_fu_1219_p1;
            trunc_ln276_reg_2053_pp0_iter1_reg <= trunc_ln276_reg_2053;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage46_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)) | ((1'b0 == ap_block_pp0_stage39_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage32_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)) | ((1'b0 == ap_block_pp0_stage25_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)) | ((1'b0 == ap_block_pp0_stage18_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            reg_1094 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage47_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)) | ((1'b0 == ap_block_pp0_stage40_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage33_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)) | ((1'b0 == ap_block_pp0_stage26_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)) | ((1'b0 == ap_block_pp0_stage19_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            reg_1100 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage48_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)) | ((1'b0 == ap_block_pp0_stage41_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)) | ((1'b0 == ap_block_pp0_stage34_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage27_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage20_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)))) begin
            reg_1106 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage49_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage42_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)) | ((1'b0 == ap_block_pp0_stage35_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage28_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage21_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)) | ((1'b0 == ap_block_pp0_stage14_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14)))) begin
            reg_1112 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage50_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage43_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage36_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage29_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)) | ((1'b0 == ap_block_pp0_stage22_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage15_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15)))) begin
            reg_1118 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage51_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)) | ((1'b0 == ap_block_pp0_stage44_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage37_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)) | ((1'b0 == ap_block_pp0_stage30_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)) | ((1'b0 == ap_block_pp0_stage23_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage16_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16)))) begin
            reg_1124 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage52_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)) | ((1'b0 == ap_block_pp0_stage45_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)) | ((1'b0 == ap_block_pp0_stage38_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage31_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)) | ((1'b0 == ap_block_pp0_stage24_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)) | ((1'b0 == ap_block_pp0_stage17_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17)))) begin
            reg_1130 <= grp_fu_1758_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage30_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)) | ((1'b0 == ap_block_pp0_stage42_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage18_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18)))) begin
            reg_1136 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage31_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)) | ((1'b0 == ap_block_pp0_stage43_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage19_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)))) begin
            reg_1142 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage44_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage20_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)) | ((1'b0 == ap_block_pp0_stage32_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)))) begin
            reg_1148 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage45_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage21_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)) | ((1'b0 == ap_block_pp0_stage33_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)))) begin
            reg_1154 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage22_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage34_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage46_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)))) begin
            reg_1159 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage23_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage35_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage47_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)))) begin
            reg_1165 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage24_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)) | ((1'b0 == ap_block_pp0_stage36_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage48_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)))) begin
            reg_1171 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage37_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)) | ((1'b0 == ap_block_pp0_stage49_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage25_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)))) begin
            reg_1177 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage38_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage50_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage26_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)))) begin
            reg_1182 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage51_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)) | ((1'b0 == ap_block_pp0_stage27_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage39_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            reg_1188 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage52_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)) | ((1'b0 == ap_block_pp0_stage28_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage40_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            reg_1194 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage29_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)) | ((1'b0 == ap_block_pp0_stage41_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            reg_1200 <= grp_fu_1754_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            this_TCurr_0_0_load_reg_2237 <= this_TCurr_0_0_q0;
            this_TCurr_0_1_load_reg_2242 <= this_TCurr_0_1_q0;
            this_TCurr_0_2_load_reg_2247 <= this_TCurr_0_2_q0;
            this_TCurr_0_3_load_reg_2252 <= this_TCurr_0_3_q0;
            this_TCurr_1_0_load_reg_2257 <= this_TCurr_1_0_q0;
            this_TCurr_1_1_load_reg_2262 <= this_TCurr_1_1_q0;
            this_TCurr_1_2_load_reg_2267 <= this_TCurr_1_2_q0;
            this_TCurr_1_3_load_reg_2272 <= this_TCurr_1_3_q0;
            this_TCurr_2_0_load_reg_2277 <= this_TCurr_2_0_q0;
            this_TCurr_2_1_load_reg_2282 <= this_TCurr_2_1_q0;
            this_TCurr_2_2_load_reg_2287 <= this_TCurr_2_2_q0;
            this_TCurr_2_3_load_reg_2292 <= this_TCurr_2_3_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            tmp_25_reg_2156 <= add_ln486_fu_1504_p2[32'd11];
            tmp_45_reg_2166 <= {{lshr_ln18_fu_1544_p2[55:53]}};
            xs_sign_reg_2146 <= data_fu_1461_p1[32'd63];
            zext_ln15_reg_2151[52 : 1] <= zext_ln15_fu_1496_p1[52 : 1];
            zext_ln18_reg_2161[31 : 0] <= zext_ln18_fu_1540_p1[31 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            tmp_301_reg_2309 <= tmp_301_fu_1996_p6;
            tmp_302_reg_2314 <= tmp_302_fu_2009_p6;
            tmp_303_reg_2319 <= tmp_303_fu_2022_p6;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            tmp_reg_2297 <= tmp_fu_1617_p3;
            val_reg_2171 <= val_fu_1574_p3;
        end
    end

    always @(*) begin
        if (((icmp_ln276_reg_2049 == 1'd1) & (1'b0 == ap_block_pp0_stage52_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
            ap_condition_exit_pp0_iter0_stage52 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage52 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage11_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11) & (icmp_ln276_reg_2049_pp0_iter1_reg == 1'd1))) begin
            ap_condition_exit_pp0_iter1_stage11 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter1_stage11 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage11_subdone) & (ap_loop_exit_ready_pp0_iter1_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b0)) begin
            ap_idle_pp0_0to0 = 1'b1;
        end else begin
            ap_idle_pp0_0to0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to2 = 1'b1;
        end else begin
            ap_idle_pp0_1to2 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage52_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            ap_sig_allocacmp_i_10 = 3'd0;
        end else begin
            ap_sig_allocacmp_i_10 = i_fu_358;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage47) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)) | ((1'b0 == ap_block_pp0_stage35) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            grp_fu_1085_p0 = reg_1200;
        end else if ((((1'b0 == ap_block_pp0_stage46) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)) | ((1'b0 == ap_block_pp0_stage34) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_1085_p0 = reg_1194;
        end else if ((((1'b0 == ap_block_pp0_stage45) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)) | ((1'b0 == ap_block_pp0_stage33) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_1085_p0 = reg_1188;
        end else if ((((1'b0 == ap_block_pp0_stage44) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage32) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_1085_p0 = reg_1182;
        end else if ((((1'b0 == ap_block_pp0_stage43) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage31) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_1085_p0 = reg_1177;
        end else if ((((1'b0 == ap_block_pp0_stage42) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)) | ((1'b0 == ap_block_pp0_stage30) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_1085_p0 = reg_1171;
        end else if ((((1'b0 == ap_block_pp0_stage41) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)) | ((1'b0 == ap_block_pp0_stage29) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_1085_p0 = reg_1165;
        end else if ((((1'b0 == ap_block_pp0_stage40) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage28) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage52) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)))) begin
            grp_fu_1085_p0 = reg_1159;
        end else if ((((1'b0 == ap_block_pp0_stage39) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage27) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage51) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)))) begin
            grp_fu_1085_p0 = reg_1154;
        end else if ((((1'b0 == ap_block_pp0_stage50) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage38) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage26) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)))) begin
            grp_fu_1085_p0 = reg_1148;
        end else if ((((1'b0 == ap_block_pp0_stage49) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage37) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)) | ((1'b0 == ap_block_pp0_stage25) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)))) begin
            grp_fu_1085_p0 = reg_1142;
        end else if ((((1'b0 == ap_block_pp0_stage48) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)) | ((1'b0 == ap_block_pp0_stage36) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage24) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)))) begin
            grp_fu_1085_p0 = reg_1136;
        end else if (((1'b0 == ap_block_pp0_stage18) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18))) begin
            grp_fu_1085_p0 = reg_1130;
        end else if (((1'b0 == ap_block_pp0_stage17) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17))) begin
            grp_fu_1085_p0 = reg_1124;
        end else if ((((1'b0 == ap_block_pp0_stage23) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage16) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16)))) begin
            grp_fu_1085_p0 = reg_1118;
        end else if ((((1'b0 == ap_block_pp0_stage22) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage15) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15)))) begin
            grp_fu_1085_p0 = reg_1112;
        end else if ((((1'b0 == ap_block_pp0_stage21) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)) | ((1'b0 == ap_block_pp0_stage14) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14)))) begin
            grp_fu_1085_p0 = reg_1106;
        end else if ((((1'b0 == ap_block_pp0_stage20) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)))) begin
            grp_fu_1085_p0 = reg_1100;
        end else if ((((1'b0 == ap_block_pp0_stage19) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            grp_fu_1085_p0 = reg_1094;
        end else begin
            grp_fu_1085_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage44) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage37) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)) | ((1'b0 == ap_block_pp0_stage30) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage51) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)))) begin
            grp_fu_1085_p1 = reg_1118;
        end else if ((((1'b0 == ap_block_pp0_stage50) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage43) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage36) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage29) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            grp_fu_1085_p1 = reg_1112;
        end else if ((((1'b0 == ap_block_pp0_stage49) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage42) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)) | ((1'b0 == ap_block_pp0_stage35) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage28) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_1085_p1 = reg_1106;
        end else if ((((1'b0 == ap_block_pp0_stage48) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)) | ((1'b0 == ap_block_pp0_stage41) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)) | ((1'b0 == ap_block_pp0_stage34) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage27) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_1085_p1 = reg_1100;
        end else if ((((1'b0 == ap_block_pp0_stage47) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)) | ((1'b0 == ap_block_pp0_stage40) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage33) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)) | ((1'b0 == ap_block_pp0_stage26) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_1085_p1 = reg_1094;
        end else if ((((1'b0 == ap_block_pp0_stage46) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)) | ((1'b0 == ap_block_pp0_stage39) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage32) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)) | ((1'b0 == ap_block_pp0_stage25) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_1085_p1 = reg_1130;
        end else if ((((1'b0 == ap_block_pp0_stage45) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)) | ((1'b0 == ap_block_pp0_stage38) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage31) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)) | ((1'b0 == ap_block_pp0_stage24) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage52) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)))) begin
            grp_fu_1085_p1 = reg_1124;
        end else if ((((1'b0 == ap_block_pp0_stage23) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage22) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage21) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)) | ((1'b0 == ap_block_pp0_stage20) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)) | ((1'b0 == ap_block_pp0_stage19) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)) | ((1'b0 == ap_block_pp0_stage18) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage17) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17)) | ((1'b0 == ap_block_pp0_stage16) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16)) | ((1'b0 == ap_block_pp0_stage15) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == 
    ap_CS_fsm_pp0_stage15)) | ((1'b0 == ap_block_pp0_stage14) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)))) begin
            grp_fu_1085_p1 = 64'd0;
        end else begin
            grp_fu_1085_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage50) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage49) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage52) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)) | ((1'b0 == ap_block_pp0_stage51) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)))) begin
            grp_fu_1090_p0 = this_TCurr_2_3_load_reg_2292;
        end else if ((((1'b0 == ap_block_pp0_stage48) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)) | ((1'b0 == ap_block_pp0_stage47) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)) | ((1'b0 == ap_block_pp0_stage46) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)) | ((1'b0 == ap_block_pp0_stage45) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)))) begin
            grp_fu_1090_p0 = this_TCurr_1_3_load_reg_2272;
        end else if ((((1'b0 == ap_block_pp0_stage44) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage43) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage42) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)) | ((1'b0 == ap_block_pp0_stage41) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)))) begin
            grp_fu_1090_p0 = this_TCurr_0_3_load_reg_2252;
        end else if ((((1'b0 == ap_block_pp0_stage40) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage39) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage38) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage37) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)))) begin
            grp_fu_1090_p0 = this_TCurr_2_2_load_reg_2287;
        end else if ((((1'b0 == ap_block_pp0_stage36) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage35) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage34) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage33) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)))) begin
            grp_fu_1090_p0 = this_TCurr_1_2_load_reg_2267;
        end else if ((((1'b0 == ap_block_pp0_stage32) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)) | ((1'b0 == ap_block_pp0_stage31) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)) | ((1'b0 == ap_block_pp0_stage30) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)) | ((1'b0 == ap_block_pp0_stage29) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)))) begin
            grp_fu_1090_p0 = this_TCurr_0_2_load_reg_2247;
        end else if ((((1'b0 == ap_block_pp0_stage28) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage27) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage26) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)) | ((1'b0 == ap_block_pp0_stage25) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)))) begin
            grp_fu_1090_p0 = this_TCurr_2_1_load_reg_2282;
        end else if ((((1'b0 == ap_block_pp0_stage24) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)) | ((1'b0 == ap_block_pp0_stage23) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage22) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage21) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)))) begin
            grp_fu_1090_p0 = this_TCurr_1_1_load_reg_2262;
        end else if ((((1'b0 == ap_block_pp0_stage20) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)) | ((1'b0 == ap_block_pp0_stage19) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)) | ((1'b0 == ap_block_pp0_stage18) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18)) | ((1'b0 == ap_block_pp0_stage17) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17)))) begin
            grp_fu_1090_p0 = this_TCurr_0_1_load_reg_2242;
        end else if ((((1'b0 == ap_block_pp0_stage16) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16)) | ((1'b0 == ap_block_pp0_stage15) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15)) | ((1'b0 == ap_block_pp0_stage14) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)))) begin
            grp_fu_1090_p0 = this_TCurr_2_0_load_reg_2277;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)))) begin
            grp_fu_1090_p0 = this_TCurr_1_0_load_reg_2257;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_1090_p0 = this_TCurr_0_0_load_reg_2237;
        end else begin
            grp_fu_1090_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage48) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage48)) | ((1'b0 == ap_block_pp0_stage44) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage44)) | ((1'b0 == ap_block_pp0_stage52) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage52)))) begin
            grp_fu_1090_p1 = tmp_300_reg_2141;
        end else if ((((1'b0 == ap_block_pp0_stage47) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage47)) | ((1'b0 == ap_block_pp0_stage43) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage43)) | ((1'b0 == ap_block_pp0_stage51) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage51)))) begin
            grp_fu_1090_p1 = tmp_296_reg_2121;
        end else if ((((1'b0 == ap_block_pp0_stage50) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage50)) | ((1'b0 == ap_block_pp0_stage46) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage46)) | ((1'b0 == ap_block_pp0_stage42) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage42)))) begin
            grp_fu_1090_p1 = tmp_292_reg_2101;
        end else if ((((1'b0 == ap_block_pp0_stage49) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage49)) | ((1'b0 == ap_block_pp0_stage45) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage45)) | ((1'b0 == ap_block_pp0_stage41) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage41)))) begin
            grp_fu_1090_p1 = tmp_288_reg_2081;
        end else if ((((1'b0 == ap_block_pp0_stage40) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage40)) | ((1'b0 == ap_block_pp0_stage36) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage36)) | ((1'b0 == ap_block_pp0_stage32) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage32)))) begin
            grp_fu_1090_p1 = tmp_299_reg_2136;
        end else if ((((1'b0 == ap_block_pp0_stage39) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage39)) | ((1'b0 == ap_block_pp0_stage35) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage35)) | ((1'b0 == ap_block_pp0_stage31) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage31)))) begin
            grp_fu_1090_p1 = tmp_295_reg_2116;
        end else if ((((1'b0 == ap_block_pp0_stage38) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage38)) | ((1'b0 == ap_block_pp0_stage34) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage34)) | ((1'b0 == ap_block_pp0_stage30) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage30)))) begin
            grp_fu_1090_p1 = tmp_291_reg_2096;
        end else if ((((1'b0 == ap_block_pp0_stage37) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage37)) | ((1'b0 == ap_block_pp0_stage33) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage33)) | ((1'b0 == ap_block_pp0_stage29) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage29)))) begin
            grp_fu_1090_p1 = tmp_287_reg_2076;
        end else if ((((1'b0 == ap_block_pp0_stage28) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage28)) | ((1'b0 == ap_block_pp0_stage24) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage24)) | ((1'b0 == ap_block_pp0_stage20) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage20)))) begin
            grp_fu_1090_p1 = tmp_298_reg_2131;
        end else if ((((1'b0 == ap_block_pp0_stage27) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage27)) | ((1'b0 == ap_block_pp0_stage23) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage23)) | ((1'b0 == ap_block_pp0_stage19) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage19)))) begin
            grp_fu_1090_p1 = tmp_294_reg_2111;
        end else if ((((1'b0 == ap_block_pp0_stage26) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage26)) | ((1'b0 == ap_block_pp0_stage22) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage22)) | ((1'b0 == ap_block_pp0_stage18) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage18)))) begin
            grp_fu_1090_p1 = tmp_290_reg_2091;
        end else if ((((1'b0 == ap_block_pp0_stage25) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage25)) | ((1'b0 == ap_block_pp0_stage21) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage21)) | ((1'b0 == ap_block_pp0_stage17) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage17)))) begin
            grp_fu_1090_p1 = tmp_286_reg_2071;
        end else if ((((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage16) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage16)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            grp_fu_1090_p1 = tmp_297_reg_2126;
        end else if ((((1'b0 == ap_block_pp0_stage15) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage15)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            grp_fu_1090_p1 = tmp_293_reg_2106;
        end else if ((((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage14) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage14)))) begin
            grp_fu_1090_p1 = tmp_289_reg_2086;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)))) begin
            grp_fu_1090_p1 = tmp_s_reg_2066;
        end else begin
            grp_fu_1090_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_0_0_constprop_o = reg_1136;
        end else begin
            l_TColl_0_0_0_constprop_o = l_TColl_0_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_0_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_0_1_constprop_o = reg_1136;
        end else begin
            l_TColl_0_0_1_constprop_o = l_TColl_0_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_0_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_0_2_constprop_o = reg_1136;
        end else begin
            l_TColl_0_0_2_constprop_o = l_TColl_0_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_0_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_0_3_constprop_o = reg_1136;
        end else begin
            l_TColl_0_0_3_constprop_o = l_TColl_0_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_0_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_1_0_constprop_o = reg_1142;
        end else begin
            l_TColl_0_1_0_constprop_o = l_TColl_0_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_1_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_1_1_constprop_o = reg_1142;
        end else begin
            l_TColl_0_1_1_constprop_o = l_TColl_0_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_1_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_1_2_constprop_o = reg_1142;
        end else begin
            l_TColl_0_1_2_constprop_o = l_TColl_0_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_1_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_1_3_constprop_o = reg_1142;
        end else begin
            l_TColl_0_1_3_constprop_o = l_TColl_0_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_1_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_2_0_constprop_o = reg_1148;
        end else begin
            l_TColl_0_2_0_constprop_o = l_TColl_0_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_2_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_2_1_constprop_o = reg_1148;
        end else begin
            l_TColl_0_2_1_constprop_o = l_TColl_0_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_2_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_2_2_constprop_o = reg_1148;
        end else begin
            l_TColl_0_2_2_constprop_o = l_TColl_0_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_2_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_2_3_constprop_o = reg_1148;
        end else begin
            l_TColl_0_2_3_constprop_o = l_TColl_0_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_2_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_3_0_constprop_o = reg_1154;
        end else begin
            l_TColl_0_3_0_constprop_o = l_TColl_0_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_0_3_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_3_1_constprop_o = reg_1154;
        end else begin
            l_TColl_0_3_1_constprop_o = l_TColl_0_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_0_3_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_3_2_constprop_o = reg_1154;
        end else begin
            l_TColl_0_3_2_constprop_o = l_TColl_0_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_0_3_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_3_3_constprop_o = reg_1154;
        end else begin
            l_TColl_0_3_3_constprop_o = l_TColl_0_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_0_3_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_0_0_constprop_o = reg_1159;
        end else begin
            l_TColl_1_0_0_constprop_o = l_TColl_1_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_0_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_0_1_constprop_o = reg_1159;
        end else begin
            l_TColl_1_0_1_constprop_o = l_TColl_1_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_0_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_0_2_constprop_o = reg_1159;
        end else begin
            l_TColl_1_0_2_constprop_o = l_TColl_1_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_0_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_0_3_constprop_o = reg_1159;
        end else begin
            l_TColl_1_0_3_constprop_o = l_TColl_1_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_0_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_1_0_constprop_o = reg_1165;
        end else begin
            l_TColl_1_1_0_constprop_o = l_TColl_1_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_1_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_1_1_constprop_o = reg_1165;
        end else begin
            l_TColl_1_1_1_constprop_o = l_TColl_1_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_1_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_1_2_constprop_o = reg_1165;
        end else begin
            l_TColl_1_1_2_constprop_o = l_TColl_1_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_1_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_1_3_constprop_o = reg_1165;
        end else begin
            l_TColl_1_1_3_constprop_o = l_TColl_1_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_1_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_2_0_constprop_o = reg_1171;
        end else begin
            l_TColl_1_2_0_constprop_o = l_TColl_1_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_2_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_2_1_constprop_o = reg_1171;
        end else begin
            l_TColl_1_2_1_constprop_o = l_TColl_1_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_2_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_2_2_constprop_o = reg_1171;
        end else begin
            l_TColl_1_2_2_constprop_o = l_TColl_1_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_2_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_2_3_constprop_o = reg_1171;
        end else begin
            l_TColl_1_2_3_constprop_o = l_TColl_1_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_2_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_3_0_constprop_o = reg_1177;
        end else begin
            l_TColl_1_3_0_constprop_o = l_TColl_1_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_1_3_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_3_1_constprop_o = reg_1177;
        end else begin
            l_TColl_1_3_1_constprop_o = l_TColl_1_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_1_3_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_3_2_constprop_o = reg_1177;
        end else begin
            l_TColl_1_3_2_constprop_o = l_TColl_1_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_1_3_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_3_3_constprop_o = reg_1177;
        end else begin
            l_TColl_1_3_3_constprop_o = l_TColl_1_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_1_3_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_0_0_constprop_o = reg_1182;
        end else begin
            l_TColl_2_0_0_constprop_o = l_TColl_2_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_0_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_0_1_constprop_o = reg_1182;
        end else begin
            l_TColl_2_0_1_constprop_o = l_TColl_2_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_0_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_0_2_constprop_o = reg_1182;
        end else begin
            l_TColl_2_0_2_constprop_o = l_TColl_2_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_0_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_0_3_constprop_o = reg_1182;
        end else begin
            l_TColl_2_0_3_constprop_o = l_TColl_2_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_0_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_1_0_constprop_o = reg_1188;
        end else begin
            l_TColl_2_1_0_constprop_o = l_TColl_2_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_1_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_1_1_constprop_o = reg_1188;
        end else begin
            l_TColl_2_1_1_constprop_o = l_TColl_2_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_1_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_1_2_constprop_o = reg_1188;
        end else begin
            l_TColl_2_1_2_constprop_o = l_TColl_2_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_1_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_1_3_constprop_o = reg_1188;
        end else begin
            l_TColl_2_1_3_constprop_o = l_TColl_2_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_1_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_2_0_constprop_o = reg_1194;
        end else begin
            l_TColl_2_2_0_constprop_o = l_TColl_2_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_2_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_2_1_constprop_o = reg_1194;
        end else begin
            l_TColl_2_2_1_constprop_o = l_TColl_2_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_2_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_2_2_constprop_o = reg_1194;
        end else begin
            l_TColl_2_2_2_constprop_o = l_TColl_2_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_2_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_2_3_constprop_o = reg_1194;
        end else begin
            l_TColl_2_2_3_constprop_o = l_TColl_2_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_2_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_3_0_constprop_o = grp_fu_1754_p_dout0;
        end else begin
            l_TColl_2_3_0_constprop_o = l_TColl_2_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd0))) begin
            l_TColl_2_3_0_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_0_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_3_1_constprop_o = grp_fu_1754_p_dout0;
        end else begin
            l_TColl_2_3_1_constprop_o = l_TColl_2_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd1))) begin
            l_TColl_2_3_1_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_1_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_3_2_constprop_o = grp_fu_1754_p_dout0;
        end else begin
            l_TColl_2_3_2_constprop_o = l_TColl_2_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd2))) begin
            l_TColl_2_3_2_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_2_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_3_3_constprop_o = grp_fu_1754_p_dout0;
        end else begin
            l_TColl_2_3_3_constprop_o = l_TColl_2_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12) & (trunc_ln276_reg_2053_pp0_iter1_reg == 2'd3))) begin
            l_TColl_2_3_3_constprop_o_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_3_constprop_o_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_0_0_ce0 = 1'b1;
        end else begin
            this_TCurr_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_0_1_ce0 = 1'b1;
        end else begin
            this_TCurr_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_0_2_ce0 = 1'b1;
        end else begin
            this_TCurr_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_0_3_ce0 = 1'b1;
        end else begin
            this_TCurr_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_1_0_ce0 = 1'b1;
        end else begin
            this_TCurr_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_1_1_ce0 = 1'b1;
        end else begin
            this_TCurr_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_1_2_ce0 = 1'b1;
        end else begin
            this_TCurr_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_1_3_ce0 = 1'b1;
        end else begin
            this_TCurr_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_2_0_ce0 = 1'b1;
        end else begin
            this_TCurr_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_2_1_ce0 = 1'b1;
        end else begin
            this_TCurr_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_2_2_ce0 = 1'b1;
        end else begin
            this_TCurr_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            this_TCurr_2_3_ce0 = 1'b1;
        end else begin
            this_TCurr_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                this_cAxes_address0 = zext_ln282_8_fu_1703_p1;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                this_cAxes_address0 = zext_ln282_5_fu_1693_p1;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                this_cAxes_address0 = zext_ln282_2_fu_1683_p1;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                this_cAxes_address0 = zext_ln282_7_fu_1673_p1;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                this_cAxes_address0 = zext_ln282_4_fu_1663_p1;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                this_cAxes_address0 = zext_ln282_1_fu_1653_p1;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                this_cAxes_address0 = zext_ln282_6_fu_1643_p1;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                this_cAxes_address0 = zext_ln282_3_fu_1633_p1;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                this_cAxes_address0 = zext_ln282_fu_1623_p1;
            end else begin
                this_cAxes_address0 = 'bx;
            end
        end else begin
            this_cAxes_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            this_cAxes_ce0 = 1'b1;
        end else begin
            this_cAxes_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                this_cAxes_d0 = reg_1194;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                this_cAxes_d0 = reg_1188;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                this_cAxes_d0 = reg_1182;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                this_cAxes_d0 = reg_1171;
            end else if (((1'b0 == ap_block_pp0_stage7) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                this_cAxes_d0 = reg_1165;
            end else if (((1'b0 == ap_block_pp0_stage6) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                this_cAxes_d0 = reg_1159;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                this_cAxes_d0 = reg_1148;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                this_cAxes_d0 = reg_1142;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                this_cAxes_d0 = reg_1136;
            end else begin
                this_cAxes_d0 = 'bx;
            end
        end else begin
            this_cAxes_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            this_cAxes_we0 = 1'b1;
        end else begin
            this_cAxes_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to2 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if (((ap_idle_pp0_0to0 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter1_stage11))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            ap_ST_fsm_pp0_stage14: begin
                if ((1'b0 == ap_block_pp0_stage14_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end
            end
            ap_ST_fsm_pp0_stage15: begin
                if ((1'b0 == ap_block_pp0_stage15_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end
            end
            ap_ST_fsm_pp0_stage16: begin
                if ((1'b0 == ap_block_pp0_stage16_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end
            end
            ap_ST_fsm_pp0_stage17: begin
                if ((1'b0 == ap_block_pp0_stage17_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end
            end
            ap_ST_fsm_pp0_stage18: begin
                if ((1'b0 == ap_block_pp0_stage18_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end
            end
            ap_ST_fsm_pp0_stage19: begin
                if ((1'b0 == ap_block_pp0_stage19_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end
            end
            ap_ST_fsm_pp0_stage20: begin
                if ((1'b0 == ap_block_pp0_stage20_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end
            end
            ap_ST_fsm_pp0_stage21: begin
                if ((1'b0 == ap_block_pp0_stage21_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end
            end
            ap_ST_fsm_pp0_stage22: begin
                if ((1'b0 == ap_block_pp0_stage22_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end
            end
            ap_ST_fsm_pp0_stage23: begin
                if ((1'b0 == ap_block_pp0_stage23_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end
            end
            ap_ST_fsm_pp0_stage24: begin
                if ((1'b0 == ap_block_pp0_stage24_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end
            end
            ap_ST_fsm_pp0_stage25: begin
                if ((1'b0 == ap_block_pp0_stage25_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end
            end
            ap_ST_fsm_pp0_stage26: begin
                if ((1'b0 == ap_block_pp0_stage26_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end
            end
            ap_ST_fsm_pp0_stage27: begin
                if ((1'b0 == ap_block_pp0_stage27_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end
            end
            ap_ST_fsm_pp0_stage28: begin
                if ((1'b0 == ap_block_pp0_stage28_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end
            end
            ap_ST_fsm_pp0_stage29: begin
                if ((1'b0 == ap_block_pp0_stage29_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end
            end
            ap_ST_fsm_pp0_stage30: begin
                if ((1'b0 == ap_block_pp0_stage30_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end
            end
            ap_ST_fsm_pp0_stage31: begin
                if ((1'b0 == ap_block_pp0_stage31_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end
            end
            ap_ST_fsm_pp0_stage32: begin
                if ((1'b0 == ap_block_pp0_stage32_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end
            end
            ap_ST_fsm_pp0_stage33: begin
                if ((1'b0 == ap_block_pp0_stage33_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end
            end
            ap_ST_fsm_pp0_stage34: begin
                if ((1'b0 == ap_block_pp0_stage34_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end
            end
            ap_ST_fsm_pp0_stage35: begin
                if ((1'b0 == ap_block_pp0_stage35_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end
            end
            ap_ST_fsm_pp0_stage36: begin
                if ((1'b0 == ap_block_pp0_stage36_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end
            end
            ap_ST_fsm_pp0_stage37: begin
                if ((1'b0 == ap_block_pp0_stage37_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end
            end
            ap_ST_fsm_pp0_stage38: begin
                if ((1'b0 == ap_block_pp0_stage38_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end
            end
            ap_ST_fsm_pp0_stage39: begin
                if ((1'b0 == ap_block_pp0_stage39_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end
            end
            ap_ST_fsm_pp0_stage40: begin
                if ((1'b0 == ap_block_pp0_stage40_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end
            end
            ap_ST_fsm_pp0_stage41: begin
                if ((1'b0 == ap_block_pp0_stage41_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end
            end
            ap_ST_fsm_pp0_stage42: begin
                if ((1'b0 == ap_block_pp0_stage42_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end
            end
            ap_ST_fsm_pp0_stage43: begin
                if ((1'b0 == ap_block_pp0_stage43_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end
            end
            ap_ST_fsm_pp0_stage44: begin
                if ((1'b0 == ap_block_pp0_stage44_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end
            end
            ap_ST_fsm_pp0_stage45: begin
                if ((1'b0 == ap_block_pp0_stage45_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end
            end
            ap_ST_fsm_pp0_stage46: begin
                if ((1'b0 == ap_block_pp0_stage46_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end
            end
            ap_ST_fsm_pp0_stage47: begin
                if ((1'b0 == ap_block_pp0_stage47_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end
            end
            ap_ST_fsm_pp0_stage48: begin
                if ((1'b0 == ap_block_pp0_stage48_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end
            end
            ap_ST_fsm_pp0_stage49: begin
                if ((1'b0 == ap_block_pp0_stage49_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end
            end
            ap_ST_fsm_pp0_stage50: begin
                if ((1'b0 == ap_block_pp0_stage50_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end
            end
            ap_ST_fsm_pp0_stage51: begin
                if ((1'b0 == ap_block_pp0_stage51_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end
            end
            ap_ST_fsm_pp0_stage52: begin
                if ((1'b0 == ap_block_pp0_stage52_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln276_fu_1607_p2 = (i_10_reg_2042 + 3'd1);

    assign add_ln282_1_fu_1678_p2 = (tmp_reg_2297 + 6'd2);

    assign add_ln282_2_fu_1628_p2 = (tmp_reg_2297 + 6'd3);

    assign add_ln282_3_fu_1658_p2 = (tmp_reg_2297 + 6'd4);

    assign add_ln282_4_fu_1688_p2 = (tmp_reg_2297 + 6'd5);

    assign add_ln282_5_fu_1638_p2 = (tmp_reg_2297 + 6'd6);

    assign add_ln282_6_fu_1668_p2 = (tmp_reg_2297 + 6'd7);

    assign add_ln282_7_fu_1698_p2 = (tmp_reg_2297 + 6'd8);

    assign add_ln282_fu_1648_p2 = (tmp_reg_2297 + 6'd1);

    assign add_ln486_fu_1504_p2 = ($signed(zext_ln486_fu_1500_p1) + $signed(12'd3073));

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage14 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_pp0_stage15 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_pp0_stage16 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_pp0_stage17 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_pp0_stage18 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_pp0_stage19 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage20 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_pp0_stage21 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_pp0_stage22 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_pp0_stage23 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_pp0_stage24 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_pp0_stage25 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_pp0_stage26 = ap_CS_fsm[32'd26];

    assign ap_CS_fsm_pp0_stage27 = ap_CS_fsm[32'd27];

    assign ap_CS_fsm_pp0_stage28 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_pp0_stage29 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage30 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_pp0_stage31 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_pp0_stage32 = ap_CS_fsm[32'd32];

    assign ap_CS_fsm_pp0_stage33 = ap_CS_fsm[32'd33];

    assign ap_CS_fsm_pp0_stage34 = ap_CS_fsm[32'd34];

    assign ap_CS_fsm_pp0_stage35 = ap_CS_fsm[32'd35];

    assign ap_CS_fsm_pp0_stage36 = ap_CS_fsm[32'd36];

    assign ap_CS_fsm_pp0_stage37 = ap_CS_fsm[32'd37];

    assign ap_CS_fsm_pp0_stage38 = ap_CS_fsm[32'd38];

    assign ap_CS_fsm_pp0_stage39 = ap_CS_fsm[32'd39];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage40 = ap_CS_fsm[32'd40];

    assign ap_CS_fsm_pp0_stage41 = ap_CS_fsm[32'd41];

    assign ap_CS_fsm_pp0_stage42 = ap_CS_fsm[32'd42];

    assign ap_CS_fsm_pp0_stage43 = ap_CS_fsm[32'd43];

    assign ap_CS_fsm_pp0_stage44 = ap_CS_fsm[32'd44];

    assign ap_CS_fsm_pp0_stage45 = ap_CS_fsm[32'd45];

    assign ap_CS_fsm_pp0_stage46 = ap_CS_fsm[32'd46];

    assign ap_CS_fsm_pp0_stage47 = ap_CS_fsm[32'd47];

    assign ap_CS_fsm_pp0_stage48 = ap_CS_fsm[32'd48];

    assign ap_CS_fsm_pp0_stage49 = ap_CS_fsm[32'd49];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage50 = ap_CS_fsm[32'd50];

    assign ap_CS_fsm_pp0_stage51 = ap_CS_fsm[32'd51];

    assign ap_CS_fsm_pp0_stage52 = ap_CS_fsm[32'd52];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage52;

    assign data_fu_1461_p1 = dc_reg_2061;

    assign grp_blockDescToBoundingBox_double_s_fu_979_ap_start = grp_blockDescToBoundingBox_double_s_fu_979_ap_start_reg;

    assign grp_fu_1754_p_ce = 1'b1;

    assign grp_fu_1754_p_din0 = grp_fu_1085_p0;

    assign grp_fu_1754_p_din1 = grp_fu_1085_p1;

    assign grp_fu_1754_p_opcode = 2'd0;

    assign grp_fu_1758_p_ce = 1'b1;

    assign grp_fu_1758_p_din0 = grp_fu_1090_p0;

    assign grp_fu_1758_p_din1 = grp_fu_1090_p1;

    assign icmp_ln276_fu_1213_p2 = ((ap_sig_allocacmp_i_10 == 3'd4) ? 1'b1 : 1'b0);

    assign lshr_ln18_fu_1544_p2 = zext_ln15_fu_1496_p1 >> zext_ln18_fu_1540_p1;

    assign mantissa_fu_1486_p4 = {{{{1'd1}, {trunc_ln505_fu_1482_p1}}}, {1'd0}};

    assign result_2_fu_1580_p2 = (3'd0 - val_reg_2171);

    assign result_fu_1585_p3 = ((xs_sign_reg_2146[0:0] == 1'b1) ? result_2_fu_1580_p2 : val_reg_2171);

    assign select_ln18_fu_1528_p3 = ((tmp_25_fu_1510_p3[0:0] == 1'b1) ? sext_ln18_fu_1524_p1 : add_ln486_fu_1504_p2);

    assign sext_ln18_1_fu_1536_p1 = $signed(select_ln18_fu_1528_p3);

    assign sext_ln18_fu_1524_p1 = $signed(sub_ln18_fu_1518_p2);

    assign shl_ln18_fu_1560_p2 = zext_ln15_reg_2151 << zext_ln18_reg_2161;

    assign sub_ln18_fu_1518_p2 = (11'd1023 - xs_exp_fu_1472_p4);

    assign this_TCurr_0_0_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_0_1_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_0_2_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_0_3_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_1_0_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_1_1_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_1_2_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_1_3_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_2_0_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_2_1_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_2_2_address0 = zext_ln278_fu_1591_p1;

    assign this_TCurr_2_3_address0 = zext_ln278_fu_1591_p1;

    assign this_cPoints_address0 = grp_blockDescToBoundingBox_double_s_fu_979_corners_address0;

    assign this_cPoints_address1 = grp_blockDescToBoundingBox_double_s_fu_979_corners_address1;

    assign this_cPoints_ce0 = grp_blockDescToBoundingBox_double_s_fu_979_corners_ce0;

    assign this_cPoints_ce1 = grp_blockDescToBoundingBox_double_s_fu_979_corners_ce1;

    assign this_cPoints_d0 = grp_blockDescToBoundingBox_double_s_fu_979_corners_d0;

    assign this_cPoints_d1 = grp_blockDescToBoundingBox_double_s_fu_979_corners_d1;

    assign this_cPoints_we0 = grp_blockDescToBoundingBox_double_s_fu_979_corners_we0;

    assign this_cPoints_we1 = grp_blockDescToBoundingBox_double_s_fu_979_corners_we1;

    assign tmp_25_fu_1510_p3 = add_ln486_fu_1504_p2[32'd11];

    assign tmp_46_fu_1564_p4 = {{shl_ln18_fu_1560_p2[55:53]}};

    assign tmp_fu_1617_p3 = {{i_10_reg_2042_pp0_iter1_reg}, {i_10_reg_2042_pp0_iter1_reg}};

    assign trunc_ln276_fu_1219_p1 = ap_sig_allocacmp_i_10[1:0];

    assign trunc_ln505_fu_1482_p1 = data_fu_1461_p1[51:0];

    assign val_fu_1574_p3 = ((tmp_25_reg_2156[0:0] == 1'b1) ? tmp_45_reg_2166 : tmp_46_fu_1564_p4);

    assign xs_exp_fu_1472_p4 = {{data_fu_1461_p1[62:52]}};

    assign zext_ln15_fu_1496_p1 = mantissa_fu_1486_p4;

    assign zext_ln18_fu_1540_p1 = $unsigned(sext_ln18_1_fu_1536_p1);

    assign zext_ln278_fu_1591_p1 = result_fu_1585_p3;

    assign zext_ln282_1_fu_1653_p1 = add_ln282_fu_1648_p2;

    assign zext_ln282_2_fu_1683_p1 = add_ln282_1_fu_1678_p2;

    assign zext_ln282_3_fu_1633_p1 = add_ln282_2_fu_1628_p2;

    assign zext_ln282_4_fu_1663_p1 = add_ln282_3_fu_1658_p2;

    assign zext_ln282_5_fu_1693_p1 = add_ln282_4_fu_1688_p2;

    assign zext_ln282_6_fu_1643_p1 = add_ln282_5_fu_1638_p2;

    assign zext_ln282_7_fu_1673_p1 = add_ln282_6_fu_1668_p2;

    assign zext_ln282_8_fu_1703_p1 = add_ln282_7_fu_1698_p2;

    assign zext_ln282_fu_1623_p1 = tmp_fu_1617_p3;

    assign zext_ln486_fu_1500_p1 = xs_exp_fu_1472_p4;

    always @(posedge ap_clk) begin
        zext_ln15_reg_2151[0] <= 1'b0;
        zext_ln15_reg_2151[136:53] <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        zext_ln18_reg_2161[136:32] <= 105'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_detectCollNode_Pipeline_VITIS_LOOP_276_1
