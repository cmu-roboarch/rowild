/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_invert4x4Matrix_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    m_address0,
    m_ce0,
    m_q0,
    m_address1,
    m_ce1,
    m_q1,
    invOut_address0,
    invOut_ce0,
    invOut_we0,
    invOut_d0
);

    parameter ap_ST_fsm_state1 = 17'd1;
    parameter ap_ST_fsm_state2 = 17'd2;
    parameter ap_ST_fsm_state3 = 17'd4;
    parameter ap_ST_fsm_state4 = 17'd8;
    parameter ap_ST_fsm_state5 = 17'd16;
    parameter ap_ST_fsm_state6 = 17'd32;
    parameter ap_ST_fsm_state7 = 17'd64;
    parameter ap_ST_fsm_state8 = 17'd128;
    parameter ap_ST_fsm_state9 = 17'd256;
    parameter ap_ST_fsm_state10 = 17'd512;
    parameter ap_ST_fsm_state11 = 17'd1024;
    parameter ap_ST_fsm_state12 = 17'd2048;
    parameter ap_ST_fsm_state13 = 17'd4096;
    parameter ap_ST_fsm_state14 = 17'd8192;
    parameter ap_ST_fsm_state15 = 17'd16384;
    parameter ap_ST_fsm_state16 = 17'd32768;
    parameter ap_ST_fsm_state17 = 17'd65536;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [3:0] m_address0;
    output m_ce0;
    input [63:0] m_q0;
    output [3:0] m_address1;
    output m_ce1;
    input [63:0] m_q1;
    output [3:0] invOut_address0;
    output invOut_ce0;
    output invOut_we0;
    output [63:0] invOut_d0;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg [3:0] m_address0;
    reg m_ce0;
    reg [3:0] m_address1;
    reg m_ce1;

    (* fsm_encoding = "none" *) reg [16:0] ap_CS_fsm;
    wire ap_CS_fsm_state1;
    wire [63:0] grp_fu_388_p2;
    reg [63:0] reg_1033;
    wire ap_CS_fsm_state7;
    wire ap_CS_fsm_state9;
    wire [63:0] grp_fu_402_p2;
    reg [63:0] reg_1039;
    wire ap_CS_fsm_state10;
    wire [63:0] grp_fu_384_p2;
    reg [63:0] reg_1046;
    wire ap_CS_fsm_state8;
    wire [63:0] grp_fu_393_p2;
    reg [63:0] reg_1052;
    wire [63:0] grp_fu_641_p2;
    reg [63:0] reg_1058;
    wire [63:0] grp_fu_420_p2;
    reg [63:0] reg_1068;
    wire ap_CS_fsm_state2;
    reg [63:0] m_load_reg_1200;
    reg [63:0] m_load_1_reg_1215;
    wire ap_CS_fsm_state3;
    reg [63:0] m_load_2_reg_1245;
    reg [63:0] m_load_3_reg_1265;
    wire ap_CS_fsm_state4;
    reg [63:0] m_load_4_reg_1292;
    reg [63:0] m_load_5_reg_1313;
    wire ap_CS_fsm_state5;
    reg [63:0] m_load_6_reg_1342;
    reg [63:0] m_load_7_reg_1358;
    wire ap_CS_fsm_state6;
    wire [63:0] grp_fu_364_p2;
    reg [63:0] sub1_reg_1382;
    reg [63:0] m_load_8_reg_1387;
    reg [63:0] m_load_9_reg_1406;
    wire [63:0] grp_fu_369_p2;
    reg [63:0] sub2_reg_1427;
    reg [63:0] m_load_10_reg_1432;
    wire [63:0] grp_fu_379_p2;
    reg [63:0] add3_reg_1440;
    reg [63:0] m_load_11_reg_1445;
    reg [63:0] add4_reg_1465;
    reg [63:0] m_load_12_reg_1470;
    wire [63:0] grp_fu_397_p2;
    reg [63:0] add10_reg_1478;
    reg [63:0] m_load_13_reg_1483;
    wire [63:0] grp_fu_411_p2;
    reg [63:0] sub21_reg_1492;
    wire [63:0] grp_fu_614_p2;
    reg [63:0] mul57_reg_1497;
    wire [63:0] grp_fu_624_p2;
    reg [63:0] mul59_reg_1503;
    wire [63:0] grp_fu_636_p2;
    reg [63:0] mul61_reg_1509;
    wire [63:0] grp_fu_661_p2;
    reg [63:0] mul68_reg_1517;
    wire [63:0] grp_fu_701_p2;
    reg [63:0] mul71_reg_1523;
    wire [63:0] grp_fu_437_p2;
    reg [63:0] sub22_reg_1531;
    wire [63:0] sub23_fu_451_p2;
    reg [63:0] sub23_reg_1536;
    wire [63:0] add25_fu_465_p2;
    reg [63:0] add25_reg_1541;
    wire [63:0] sub28_fu_479_p2;
    reg [63:0] sub28_reg_1546;
    wire [63:0] add32_fu_493_p2;
    reg [63:0] add32_reg_1551;
    wire [63:0] add33_fu_507_p2;
    reg [63:0] add33_reg_1556;
    wire [63:0] sub35_fu_521_p2;
    reg [63:0] sub35_reg_1561;
    wire [63:0] add38_fu_535_p2;
    reg [63:0] add38_reg_1566;
    wire [63:0] det_2_fu_549_p2;
    reg [63:0] det_2_reg_1571;
    wire [63:0] grp_fu_416_p2;
    reg [63:0] add29_reg_1577;
    wire [63:0] grp_fu_428_p2;
    reg [63:0] sub34_reg_1582;
    reg [63:0] add37_reg_1587;
    wire [63:0] grp_fu_446_p2;
    reg [63:0] sub39_reg_1592;
    wire [0:0] and_ln149_fu_1174_p2;
    reg [0:0] and_ln149_reg_1597;
    wire ap_CS_fsm_state15;
    wire [63:0] grp_fu_1022_p2;
    reg [63:0] det_reg_1601;
    wire ap_CS_fsm_state16;
    reg [3:0] inv_address0;
    reg inv_ce0;
    reg inv_we0;
    reg [63:0] inv_d0;
    wire [63:0] inv_q0;
    reg [3:0] inv_address1;
    reg inv_ce1;
    reg inv_we1;
    reg [63:0] inv_d1;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_done;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_idle;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_ready;
    wire   [3:0] grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_address0;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_ce0;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_we0;
    wire   [63:0] grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_d0;
    wire   [3:0] grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_address0;
    wire grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_ce0;
    reg grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg;
    wire ap_CS_fsm_state17;
    wire ap_CS_fsm_state11;
    wire ap_CS_fsm_state12;
    wire ap_CS_fsm_state13;
    wire ap_CS_fsm_state14;
    wire [63:0] grp_fu_375_p2;
    reg [63:0] grp_fu_360_p0;
    wire [63:0] grp_fu_560_p2;
    reg [63:0] grp_fu_360_p1;
    wire [63:0] grp_fu_570_p2;
    wire [63:0] grp_fu_556_p2;
    wire [63:0] grp_fu_360_p2;
    reg [63:0] grp_fu_364_p1;
    wire [63:0] grp_fu_580_p2;
    wire [63:0] grp_fu_566_p2;
    reg [63:0] grp_fu_369_p0;
    reg [63:0] grp_fu_369_p1;
    wire [63:0] grp_fu_576_p2;
    reg [63:0] grp_fu_375_p0;
    wire [63:0] grp_fu_593_p2;
    reg [63:0] grp_fu_375_p1;
    wire [63:0] grp_fu_603_p2;
    wire [63:0] grp_fu_589_p2;
    reg [63:0] grp_fu_379_p0;
    wire [63:0] grp_fu_599_p2;
    reg [63:0] grp_fu_379_p1;
    wire [63:0] grp_fu_609_p2;
    reg [63:0] grp_fu_384_p0;
    reg [63:0] grp_fu_384_p1;
    wire [63:0] grp_fu_630_p2;
    wire [63:0] grp_fu_620_p2;
    reg [63:0] grp_fu_388_p0;
    reg [63:0] grp_fu_388_p1;
    reg [63:0] grp_fu_393_p0;
    wire [63:0] grp_fu_651_p2;
    reg [63:0] grp_fu_393_p1;
    wire [63:0] grp_fu_657_p2;
    reg [63:0] grp_fu_397_p0;
    reg [63:0] grp_fu_397_p1;
    wire [63:0] grp_fu_667_p2;
    reg [63:0] grp_fu_402_p0;
    reg [63:0] grp_fu_402_p1;
    wire [63:0] grp_fu_673_p2;
    reg [63:0] grp_fu_411_p0;
    wire [63:0] grp_fu_711_p2;
    reg [63:0] grp_fu_411_p1;
    wire [63:0] grp_fu_717_p2;
    reg [63:0] grp_fu_416_p0;
    wire [63:0] grp_fu_705_p2;
    reg [63:0] grp_fu_416_p1;
    wire [63:0] mul77_fu_751_p2;
    reg [63:0] grp_fu_420_p0;
    reg [63:0] grp_fu_420_p1;
    wire [63:0] mul78_fu_757_p2;
    reg [63:0] grp_fu_428_p0;
    reg [63:0] grp_fu_428_p1;
    wire [63:0] mul88_fu_768_p2;
    reg [63:0] grp_fu_432_p0;
    reg [63:0] grp_fu_432_p1;
    wire [63:0] mul89_fu_774_p2;
    wire [63:0] grp_fu_432_p2;
    reg [63:0] grp_fu_437_p1;
    wire [63:0] mul90_fu_780_p2;
    reg [63:0] grp_fu_442_p0;
    wire [63:0] mul92_fu_790_p2;
    reg [63:0] grp_fu_442_p1;
    wire [63:0] mul94_fu_801_p2;
    wire [63:0] grp_fu_442_p2;
    reg [63:0] grp_fu_446_p1;
    wire [63:0] mul96_fu_811_p2;
    wire [63:0] grp_fu_647_p2;
    wire [63:0] mul98_fu_822_p2;
    wire [63:0] mul102_fu_833_p2;
    wire [63:0] mul103_fu_839_p2;
    wire [63:0] sub25_fu_456_p2;
    wire [63:0] mul105_fu_849_p2;
    wire [63:0] sub26_fu_460_p2;
    wire [63:0] mul106_fu_855_p2;
    wire [63:0] mul110_fu_865_p2;
    wire [63:0] mul112_fu_876_p2;
    wire [63:0] add27_fu_470_p2;
    wire [63:0] mul113_fu_882_p2;
    wire [63:0] add28_fu_474_p2;
    wire [63:0] mul114_fu_888_p2;
    wire [63:0] mul121_fu_894_p2;
    wire [63:0] sub30_fu_484_p2;
    wire [63:0] mul122_fu_900_p2;
    wire [63:0] sub31_fu_488_p2;
    wire [63:0] mul123_fu_905_p2;
    wire [63:0] mul124_fu_911_p2;
    wire [63:0] mul125_fu_917_p2;
    wire [63:0] sub32_fu_498_p2;
    wire [63:0] mul126_fu_923_p2;
    wire [63:0] sub33_fu_502_p2;
    wire [63:0] mul127_fu_929_p2;
    wire [63:0] mul130_fu_935_p2;
    wire [63:0] mul131_fu_941_p2;
    wire [63:0] add35_fu_512_p2;
    wire [63:0] mul132_fu_947_p2;
    wire [63:0] add36_fu_516_p2;
    wire [63:0] mul133_fu_953_p2;
    wire [63:0] mul136_fu_959_p2;
    wire [63:0] mul137_fu_965_p2;
    wire [63:0] sub37_fu_526_p2;
    wire [63:0] mul138_fu_971_p2;
    wire [63:0] sub38_fu_530_p2;
    wire [63:0] mul139_fu_977_p2;
    wire [63:0] mul142_fu_983_p2;
    wire [63:0] mul143_fu_989_p2;
    wire [63:0] add40_fu_540_p2;
    wire [63:0] mul144_fu_994_p2;
    wire [63:0] add41_fu_544_p2;
    wire [63:0] mul145_fu_999_p2;
    reg [63:0] grp_fu_556_p0;
    reg [63:0] grp_fu_556_p1;
    reg [63:0] grp_fu_560_p0;
    reg [63:0] grp_fu_560_p1;
    reg [63:0] grp_fu_566_p0;
    reg [63:0] grp_fu_566_p1;
    reg [63:0] grp_fu_570_p0;
    reg [63:0] grp_fu_570_p1;
    reg [63:0] grp_fu_576_p0;
    reg [63:0] grp_fu_576_p1;
    reg [63:0] grp_fu_580_p0;
    reg [63:0] grp_fu_580_p1;
    reg [63:0] grp_fu_589_p0;
    reg [63:0] grp_fu_589_p1;
    wire [63:0] bitcast_ln42_1_fu_1083_p1;
    reg [63:0] grp_fu_593_p0;
    reg [63:0] grp_fu_593_p1;
    reg [63:0] grp_fu_599_p0;
    reg [63:0] grp_fu_599_p1;
    reg [63:0] grp_fu_603_p0;
    reg [63:0] grp_fu_603_p1;
    reg [63:0] grp_fu_609_p0;
    reg [63:0] grp_fu_609_p1;
    reg [63:0] grp_fu_614_p0;
    reg [63:0] grp_fu_614_p1;
    reg [63:0] grp_fu_620_p0;
    reg [63:0] grp_fu_620_p1;
    wire [63:0] bitcast_ln63_1_fu_1099_p1;
    reg [63:0] grp_fu_624_p0;
    reg [63:0] grp_fu_624_p1;
    reg [63:0] grp_fu_630_p0;
    reg [63:0] grp_fu_630_p1;
    reg [63:0] grp_fu_636_p0;
    reg [63:0] grp_fu_636_p1;
    reg [63:0] grp_fu_641_p0;
    reg [63:0] grp_fu_641_p1;
    reg [63:0] grp_fu_647_p0;
    reg [63:0] grp_fu_647_p1;
    wire [63:0] bitcast_ln77_1_fu_1115_p1;
    reg [63:0] grp_fu_651_p1;
    reg [63:0] grp_fu_657_p0;
    reg [63:0] grp_fu_657_p1;
    reg [63:0] grp_fu_661_p0;
    reg [63:0] grp_fu_661_p1;
    reg [63:0] grp_fu_667_p0;
    reg [63:0] grp_fu_667_p1;
    reg [63:0] grp_fu_673_p0;
    reg [63:0] grp_fu_673_p1;
    reg [63:0] grp_fu_701_p0;
    reg [63:0] grp_fu_701_p1;
    reg [63:0] grp_fu_705_p0;
    reg [63:0] grp_fu_705_p1;
    reg [63:0] grp_fu_711_p0;
    reg [63:0] grp_fu_711_p1;
    reg [63:0] grp_fu_717_p0;
    reg [63:0] grp_fu_717_p1;
    wire [63:0] mul87_fu_763_p2;
    wire [63:0] mul91_fu_786_p2;
    wire [63:0] mul93_fu_796_p2;
    wire [63:0] mul95_fu_807_p2;
    wire [63:0] mul97_fu_817_p2;
    wire [63:0] mul101_fu_828_p2;
    wire [63:0] mul104_fu_845_p2;
    wire [63:0] mul109_fu_861_p2;
    wire [63:0] mul111_fu_871_p2;
    wire [63:0] tmp_3_fu_1028_p0;
    wire [63:0] bitcast_ln42_fu_1074_p1;
    wire [63:0] xor_ln42_fu_1077_p2;
    wire [63:0] bitcast_ln63_fu_1089_p1;
    wire [63:0] xor_ln63_fu_1093_p2;
    wire [63:0] bitcast_ln77_fu_1105_p1;
    wire [63:0] xor_ln77_fu_1109_p2;
    wire [63:0] data_fu_1122_p1;
    wire [62:0] trunc_ln479_fu_1125_p1;
    wire [63:0] t_fu_1133_p3;
    wire [10:0] tmp_2_fu_1146_p4;
    wire [51:0] trunc_ln149_fu_1129_p1;
    wire [0:0] icmp_ln149_1_fu_1162_p2;
    wire [0:0] icmp_ln149_fu_1156_p2;
    wire [0:0] or_ln149_fu_1168_p2;
    wire [0:0] tmp_3_fu_1028_p2;
    reg [1:0] grp_fu_360_opcode;
    reg [1:0] grp_fu_364_opcode;
    reg [1:0] grp_fu_369_opcode;
    reg [1:0] grp_fu_379_opcode;
    reg [1:0] grp_fu_388_opcode;
    reg [1:0] grp_fu_416_opcode;
    reg [1:0] grp_fu_428_opcode;
    reg [1:0] grp_fu_432_opcode;
    reg [1:0] grp_fu_437_opcode;
    reg [1:0] grp_fu_446_opcode;
    reg ap_block_state17_on_subcall_done;
    reg [16:0] ap_NS_fsm;
    reg ap_ST_fsm_state1_blk;
    wire ap_ST_fsm_state2_blk;
    wire ap_ST_fsm_state3_blk;
    wire ap_ST_fsm_state4_blk;
    wire ap_ST_fsm_state5_blk;
    wire ap_ST_fsm_state6_blk;
    wire ap_ST_fsm_state7_blk;
    wire ap_ST_fsm_state8_blk;
    wire ap_ST_fsm_state9_blk;
    wire ap_ST_fsm_state10_blk;
    wire ap_ST_fsm_state11_blk;
    wire ap_ST_fsm_state12_blk;
    wire ap_ST_fsm_state13_blk;
    wire ap_ST_fsm_state14_blk;
    wire ap_ST_fsm_state15_blk;
    wire ap_ST_fsm_state16_blk;
    reg ap_ST_fsm_state17_blk;
    wire ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 17'd1;
        #0
        grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg = 1'b0;
    end

    main_invert4x4Matrix_double_s_inv_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(16),
        .AddressWidth(4)
    ) inv_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(inv_address0),
        .ce0(inv_ce0),
        .we0(inv_we0),
        .d0(inv_d0),
        .q0(inv_q0),
        .address1(inv_address1),
        .ce1(inv_ce1),
        .we1(inv_we1),
        .d1(inv_d1)
    );

    main_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2 grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start),
        .ap_done(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_done),
        .ap_idle(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_idle),
        .ap_ready(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_ready),
        .invOut_address0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_address0),
        .invOut_ce0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_ce0),
        .invOut_we0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_we0),
        .invOut_d0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_d0),
        .inv_address0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_address0),
        .inv_ce0(grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_ce0),
        .inv_q0(inv_q0),
        .det(det_reg_1601)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U6 (
        .din0  (grp_fu_360_p0),
        .din1  (grp_fu_360_p1),
        .opcode(grp_fu_360_opcode),
        .dout  (grp_fu_360_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U7 (
        .din0  (grp_fu_360_p2),
        .din1  (grp_fu_364_p1),
        .opcode(grp_fu_364_opcode),
        .dout  (grp_fu_364_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U8 (
        .din0  (grp_fu_369_p0),
        .din1  (grp_fu_369_p1),
        .opcode(grp_fu_369_opcode),
        .dout  (grp_fu_369_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U9 (
        .din0(grp_fu_375_p0),
        .din1(grp_fu_375_p1),
        .dout(grp_fu_375_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U10 (
        .din0  (grp_fu_379_p0),
        .din1  (grp_fu_379_p1),
        .opcode(grp_fu_379_opcode),
        .dout  (grp_fu_379_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U11 (
        .din0(grp_fu_384_p0),
        .din1(grp_fu_384_p1),
        .dout(grp_fu_384_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U12 (
        .din0  (grp_fu_388_p0),
        .din1  (grp_fu_388_p1),
        .opcode(grp_fu_388_opcode),
        .dout  (grp_fu_388_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U13 (
        .din0(grp_fu_393_p0),
        .din1(grp_fu_393_p1),
        .dout(grp_fu_393_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U14 (
        .din0(grp_fu_397_p0),
        .din1(grp_fu_397_p1),
        .dout(grp_fu_397_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U15 (
        .din0(grp_fu_402_p0),
        .din1(grp_fu_402_p1),
        .dout(grp_fu_402_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U16 (
        .din0(grp_fu_411_p0),
        .din1(grp_fu_411_p1),
        .dout(grp_fu_411_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U17 (
        .din0  (grp_fu_416_p0),
        .din1  (grp_fu_416_p1),
        .opcode(grp_fu_416_opcode),
        .dout  (grp_fu_416_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U18 (
        .din0(grp_fu_420_p0),
        .din1(grp_fu_420_p1),
        .dout(grp_fu_420_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U19 (
        .din0  (grp_fu_428_p0),
        .din1  (grp_fu_428_p1),
        .opcode(grp_fu_428_opcode),
        .dout  (grp_fu_428_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U20 (
        .din0  (grp_fu_432_p0),
        .din1  (grp_fu_432_p1),
        .opcode(grp_fu_432_opcode),
        .dout  (grp_fu_432_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U21 (
        .din0  (grp_fu_432_p2),
        .din1  (grp_fu_437_p1),
        .opcode(grp_fu_437_opcode),
        .dout  (grp_fu_437_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U22 (
        .din0(grp_fu_442_p0),
        .din1(grp_fu_442_p1),
        .dout(grp_fu_442_p2)
    );

    main_dadddsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_1_full_dsp_1_U23 (
        .din0  (grp_fu_442_p2),
        .din1  (grp_fu_446_p1),
        .opcode(grp_fu_446_opcode),
        .dout  (grp_fu_446_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U24 (
        .din0(grp_fu_446_p2),
        .din1(mul98_fu_822_p2),
        .dout(sub23_fu_451_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U25 (
        .din0(mul102_fu_833_p2),
        .din1(mul103_fu_839_p2),
        .dout(sub25_fu_456_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U26 (
        .din0(sub25_fu_456_p2),
        .din1(mul105_fu_849_p2),
        .dout(sub26_fu_460_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U27 (
        .din0(sub26_fu_460_p2),
        .din1(mul106_fu_855_p2),
        .dout(add25_fu_465_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U28 (
        .din0(mul110_fu_865_p2),
        .din1(mul112_fu_876_p2),
        .dout(add27_fu_470_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U29 (
        .din0(add27_fu_470_p2),
        .din1(mul113_fu_882_p2),
        .dout(add28_fu_474_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U30 (
        .din0(add28_fu_474_p2),
        .din1(mul114_fu_888_p2),
        .dout(sub28_fu_479_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U31 (
        .din0(reg_1068),
        .din1(mul121_fu_894_p2),
        .dout(sub30_fu_484_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U32 (
        .din0(sub30_fu_484_p2),
        .din1(mul122_fu_900_p2),
        .dout(sub31_fu_488_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U33 (
        .din0(sub31_fu_488_p2),
        .din1(mul123_fu_905_p2),
        .dout(add32_fu_493_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U34 (
        .din0(mul124_fu_911_p2),
        .din1(mul125_fu_917_p2),
        .dout(sub32_fu_498_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U35 (
        .din0(sub32_fu_498_p2),
        .din1(mul126_fu_923_p2),
        .dout(sub33_fu_502_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U36 (
        .din0(sub33_fu_502_p2),
        .din1(mul127_fu_929_p2),
        .dout(add33_fu_507_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U37 (
        .din0(mul130_fu_935_p2),
        .din1(mul131_fu_941_p2),
        .dout(add35_fu_512_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U38 (
        .din0(add35_fu_512_p2),
        .din1(mul132_fu_947_p2),
        .dout(add36_fu_516_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U39 (
        .din0(add36_fu_516_p2),
        .din1(mul133_fu_953_p2),
        .dout(sub35_fu_521_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U40 (
        .din0(mul136_fu_959_p2),
        .din1(mul137_fu_965_p2),
        .dout(sub37_fu_526_p2)
    );

    main_dsub_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsub_64ns_64ns_64_1_full_dsp_1_U41 (
        .din0(sub37_fu_526_p2),
        .din1(mul138_fu_971_p2),
        .dout(sub38_fu_530_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U42 (
        .din0(sub38_fu_530_p2),
        .din1(mul139_fu_977_p2),
        .dout(add38_fu_535_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U43 (
        .din0(mul142_fu_983_p2),
        .din1(mul143_fu_989_p2),
        .dout(add40_fu_540_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U44 (
        .din0(add40_fu_540_p2),
        .din1(mul144_fu_994_p2),
        .dout(add41_fu_544_p2)
    );

    main_dadd_64ns_64ns_64_1_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_1_full_dsp_1_U45 (
        .din0(add41_fu_544_p2),
        .din1(mul145_fu_999_p2),
        .dout(det_2_fu_549_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U46 (
        .din0(grp_fu_556_p0),
        .din1(grp_fu_556_p1),
        .dout(grp_fu_556_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U47 (
        .din0(grp_fu_560_p0),
        .din1(grp_fu_560_p1),
        .dout(grp_fu_560_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U48 (
        .din0(grp_fu_566_p0),
        .din1(grp_fu_566_p1),
        .dout(grp_fu_566_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U49 (
        .din0(grp_fu_570_p0),
        .din1(grp_fu_570_p1),
        .dout(grp_fu_570_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U50 (
        .din0(grp_fu_576_p0),
        .din1(grp_fu_576_p1),
        .dout(grp_fu_576_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U51 (
        .din0(grp_fu_580_p0),
        .din1(grp_fu_580_p1),
        .dout(grp_fu_580_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U52 (
        .din0(grp_fu_589_p0),
        .din1(grp_fu_589_p1),
        .dout(grp_fu_589_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U53 (
        .din0(grp_fu_593_p0),
        .din1(grp_fu_593_p1),
        .dout(grp_fu_593_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U54 (
        .din0(grp_fu_599_p0),
        .din1(grp_fu_599_p1),
        .dout(grp_fu_599_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U55 (
        .din0(grp_fu_603_p0),
        .din1(grp_fu_603_p1),
        .dout(grp_fu_603_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U56 (
        .din0(grp_fu_609_p0),
        .din1(grp_fu_609_p1),
        .dout(grp_fu_609_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U57 (
        .din0(grp_fu_614_p0),
        .din1(grp_fu_614_p1),
        .dout(grp_fu_614_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U58 (
        .din0(grp_fu_620_p0),
        .din1(grp_fu_620_p1),
        .dout(grp_fu_620_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U59 (
        .din0(grp_fu_624_p0),
        .din1(grp_fu_624_p1),
        .dout(grp_fu_624_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U60 (
        .din0(grp_fu_630_p0),
        .din1(grp_fu_630_p1),
        .dout(grp_fu_630_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U61 (
        .din0(grp_fu_636_p0),
        .din1(grp_fu_636_p1),
        .dout(grp_fu_636_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U62 (
        .din0(grp_fu_641_p0),
        .din1(grp_fu_641_p1),
        .dout(grp_fu_641_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U63 (
        .din0(grp_fu_647_p0),
        .din1(grp_fu_647_p1),
        .dout(grp_fu_647_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U64 (
        .din0(grp_fu_647_p2),
        .din1(grp_fu_651_p1),
        .dout(grp_fu_651_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U65 (
        .din0(grp_fu_657_p0),
        .din1(grp_fu_657_p1),
        .dout(grp_fu_657_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U66 (
        .din0(grp_fu_661_p0),
        .din1(grp_fu_661_p1),
        .dout(grp_fu_661_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U67 (
        .din0(grp_fu_667_p0),
        .din1(grp_fu_667_p1),
        .dout(grp_fu_667_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U68 (
        .din0(grp_fu_673_p0),
        .din1(grp_fu_673_p1),
        .dout(grp_fu_673_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U69 (
        .din0(grp_fu_701_p0),
        .din1(grp_fu_701_p1),
        .dout(grp_fu_701_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U70 (
        .din0(grp_fu_705_p0),
        .din1(grp_fu_705_p1),
        .dout(grp_fu_705_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U71 (
        .din0(grp_fu_711_p0),
        .din1(grp_fu_711_p1),
        .dout(grp_fu_711_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U72 (
        .din0(grp_fu_717_p0),
        .din1(grp_fu_717_p1),
        .dout(grp_fu_717_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U73 (
        .din0(grp_fu_661_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul77_fu_751_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U74 (
        .din0(grp_fu_614_p2),
        .din1(m_load_8_reg_1387),
        .dout(mul78_fu_757_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U75 (
        .din0(m_load_reg_1200),
        .din1(m_q1),
        .dout(mul87_fu_763_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U76 (
        .din0(mul87_fu_763_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul88_fu_768_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U77 (
        .din0(grp_fu_570_p2),
        .din1(m_load_7_reg_1358),
        .dout(mul89_fu_774_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U78 (
        .din0(grp_fu_580_p2),
        .din1(m_load_6_reg_1342),
        .dout(mul90_fu_780_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U79 (
        .din0(m_load_6_reg_1342),
        .din1(bitcast_ln77_1_fu_1115_p1),
        .dout(mul91_fu_786_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U80 (
        .din0(mul91_fu_786_p2),
        .din1(m_load_2_reg_1245),
        .dout(mul92_fu_790_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U81 (
        .din0(m_q0),
        .din1(m_load_7_reg_1358),
        .dout(mul93_fu_796_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U82 (
        .din0(mul93_fu_796_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul94_fu_801_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U83 (
        .din0(m_load_9_reg_1406),
        .din1(m_load_13_reg_1483),
        .dout(mul95_fu_807_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U84 (
        .din0(mul95_fu_807_p2),
        .din1(m_load_2_reg_1245),
        .dout(mul96_fu_811_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U85 (
        .din0(m_load_9_reg_1406),
        .din1(m_q1),
        .dout(mul97_fu_817_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U86 (
        .din0(mul97_fu_817_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul98_fu_822_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U87 (
        .din0(m_q0),
        .din1(m_load_reg_1200),
        .dout(mul101_fu_828_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U88 (
        .din0(mul101_fu_828_p2),
        .din1(m_load_2_reg_1245),
        .dout(mul102_fu_833_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U89 (
        .din0(mul93_fu_796_p2),
        .din1(m_load_8_reg_1387),
        .dout(mul103_fu_839_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U90 (
        .din0(m_load_9_reg_1406),
        .din1(m_load_12_reg_1470),
        .dout(mul104_fu_845_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U91 (
        .din0(mul104_fu_845_p2),
        .din1(m_load_2_reg_1245),
        .dout(mul105_fu_849_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U92 (
        .din0(mul97_fu_817_p2),
        .din1(m_load_8_reg_1387),
        .dout(mul106_fu_855_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U93 (
        .din0(m_load_reg_1200),
        .din1(bitcast_ln77_1_fu_1115_p1),
        .dout(mul109_fu_861_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U94 (
        .din0(mul109_fu_861_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul110_fu_865_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U95 (
        .din0(m_q0),
        .din1(m_load_6_reg_1342),
        .dout(mul111_fu_871_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U96 (
        .din0(mul111_fu_871_p2),
        .din1(m_load_8_reg_1387),
        .dout(mul112_fu_876_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U97 (
        .din0(mul104_fu_845_p2),
        .din1(m_load_4_reg_1292),
        .dout(mul113_fu_882_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U98 (
        .din0(mul95_fu_807_p2),
        .din1(m_load_8_reg_1387),
        .dout(mul114_fu_888_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U99 (
        .din0(mul87_fu_763_p2),
        .din1(m_load_1_reg_1215),
        .dout(mul121_fu_894_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U100 (
        .din0(reg_1058),
        .din1(m_load_7_reg_1358),
        .dout(mul122_fu_900_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U101 (
        .din0(grp_fu_560_p2),
        .din1(m_load_6_reg_1342),
        .dout(mul123_fu_905_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U102 (
        .din0(mul111_fu_871_p2),
        .din1(m_load_3_reg_1265),
        .dout(mul124_fu_911_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U103 (
        .din0(mul93_fu_796_p2),
        .din1(m_load_1_reg_1215),
        .dout(mul125_fu_917_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U104 (
        .din0(mul95_fu_807_p2),
        .din1(m_load_3_reg_1265),
        .dout(mul126_fu_923_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U105 (
        .din0(mul97_fu_817_p2),
        .din1(m_load_1_reg_1215),
        .dout(mul127_fu_929_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U106 (
        .din0(mul109_fu_861_p2),
        .din1(m_load_3_reg_1265),
        .dout(mul130_fu_935_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U107 (
        .din0(mul93_fu_796_p2),
        .din1(m_load_5_reg_1313),
        .dout(mul131_fu_941_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U108 (
        .din0(mul104_fu_845_p2),
        .din1(m_load_3_reg_1265),
        .dout(mul132_fu_947_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U109 (
        .din0(mul97_fu_817_p2),
        .din1(m_load_5_reg_1313),
        .dout(mul133_fu_953_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U110 (
        .din0(mul101_fu_828_p2),
        .din1(m_load_1_reg_1215),
        .dout(mul136_fu_959_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U111 (
        .din0(mul111_fu_871_p2),
        .din1(m_load_5_reg_1313),
        .dout(mul137_fu_965_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U112 (
        .din0(mul104_fu_845_p2),
        .din1(m_load_1_reg_1215),
        .dout(mul138_fu_971_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U113 (
        .din0(mul95_fu_807_p2),
        .din1(m_load_5_reg_1313),
        .dout(mul139_fu_977_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U114 (
        .din0(m_q0),
        .din1(sub2_reg_1427),
        .dout(mul142_fu_983_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U115 (
        .din0(m_load_12_reg_1470),
        .din1(add4_reg_1465),
        .dout(mul143_fu_989_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U116 (
        .din0(m_load_13_reg_1483),
        .din1(reg_1046),
        .dout(mul144_fu_994_p2)
    );

    main_dmul_64ns_64ns_64_1_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_1_max_dsp_1_U117 (
        .din0(m_q1),
        .din1(reg_1052),
        .dout(mul145_fu_999_p2)
    );

    main_ddiv_64ns_64ns_64_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) ddiv_64ns_64ns_64_2_no_dsp_1_U118 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd4607182418800017408),
        .din1(det_2_reg_1571),
        .ce(1'b1),
        .dout(grp_fu_1022_p2)
    );

    main_dcmp_64ns_64ns_1_1_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_1_no_dsp_1_U119 (
        .din0  (tmp_3_fu_1028_p0),
        .din1  (64'd4517329193108106637),
        .opcode(5'd4),
        .dout  (tmp_3_fu_1028_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state16)) begin
                grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg <= 1'b1;
            end else if ((grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_ready == 1'b1)) begin
                grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            add10_reg_1478 <= grp_fu_397_p2;
            add4_reg_1465 <= grp_fu_369_p2;
            m_load_12_reg_1470 <= m_q1;
            m_load_13_reg_1483 <= m_q0;
            sub21_reg_1492 <= grp_fu_411_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            add25_reg_1541 <= add25_fu_465_p2;
            add32_reg_1551 <= add32_fu_493_p2;
            add33_reg_1556 <= add33_fu_507_p2;
            add38_reg_1566 <= add38_fu_535_p2;
            det_2_reg_1571 <= det_2_fu_549_p2;
            mul57_reg_1497 <= grp_fu_614_p2;
            mul59_reg_1503 <= grp_fu_624_p2;
            mul61_reg_1509 <= grp_fu_636_p2;
            mul68_reg_1517 <= grp_fu_661_p2;
            mul71_reg_1523 <= grp_fu_701_p2;
            sub22_reg_1531 <= grp_fu_437_p2;
            sub23_reg_1536 <= sub23_fu_451_p2;
            sub28_reg_1546 <= sub28_fu_479_p2;
            sub35_reg_1561 <= sub35_fu_521_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            add29_reg_1577 <= grp_fu_416_p2;
            add37_reg_1587 <= grp_fu_437_p2;
            sub34_reg_1582 <= grp_fu_428_p2;
            sub39_reg_1592 <= grp_fu_446_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            add3_reg_1440 <= grp_fu_379_p2;
            m_load_10_reg_1432 <= m_q1;
            m_load_11_reg_1445 <= m_q0;
            sub2_reg_1427 <= grp_fu_369_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            and_ln149_reg_1597 <= and_ln149_fu_1174_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state16)) begin
            det_reg_1601 <= grp_fu_1022_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            m_load_1_reg_1215 <= m_q0;
            m_load_reg_1200   <= m_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            m_load_2_reg_1245 <= m_q1;
            m_load_3_reg_1265 <= m_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            m_load_4_reg_1292 <= m_q1;
            m_load_5_reg_1313 <= m_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            m_load_6_reg_1342 <= m_q1;
            m_load_7_reg_1358 <= m_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state6)) begin
            m_load_8_reg_1387 <= m_q1;
            m_load_9_reg_1406 <= m_q0;
            sub1_reg_1382 <= grp_fu_364_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            reg_1033 <= grp_fu_388_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            reg_1039 <= grp_fu_402_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10))) begin
            reg_1046 <= grp_fu_384_p2;
            reg_1052 <= grp_fu_393_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9))) begin
            reg_1058 <= grp_fu_641_p2;
            reg_1068 <= grp_fu_420_p2;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state17_on_subcall_done)) begin
            ap_ST_fsm_state17_blk = 1'b1;
        end else begin
            ap_ST_fsm_state17_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state2_blk = 1'b0;

    assign ap_ST_fsm_state3_blk = 1'b0;

    assign ap_ST_fsm_state4_blk = 1'b0;

    assign ap_ST_fsm_state5_blk = 1'b0;

    assign ap_ST_fsm_state6_blk = 1'b0;

    assign ap_ST_fsm_state7_blk = 1'b0;

    assign ap_ST_fsm_state8_blk = 1'b0;

    assign ap_ST_fsm_state9_blk = 1'b0;

    always @(*) begin
        if ((((1'b0 == ap_block_state17_on_subcall_done) & (1'b1 == ap_CS_fsm_state17)) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_state17_on_subcall_done) & (1'b1 == ap_CS_fsm_state17))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_360_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_360_opcode = 2'd0;
        end else begin
            grp_fu_360_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_360_p0 = reg_1033;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_360_p0 = add10_reg_1478;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_360_p0 = add3_reg_1440;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_360_p0 = sub1_reg_1382;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_360_p0 = grp_fu_560_p2;
        end else begin
            grp_fu_360_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_360_p1 = grp_fu_556_p2;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_360_p1 = grp_fu_560_p2;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_360_p1 = grp_fu_570_p2;
        end else begin
            grp_fu_360_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_364_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_364_opcode = 2'd0;
        end else begin
            grp_fu_364_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_364_p1 = grp_fu_560_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_364_p1 = grp_fu_566_p2;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_364_p1 = grp_fu_570_p2;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_364_p1 = grp_fu_580_p2;
        end else begin
            grp_fu_364_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_369_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_369_opcode = 2'd0;
        end else begin
            grp_fu_369_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_369_p0 = reg_1039;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_369_p0 = grp_fu_364_p2;
        end else begin
            grp_fu_369_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_369_p1 = grp_fu_566_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_369_p1 = grp_fu_576_p2;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_369_p1 = grp_fu_580_p2;
        end else begin
            grp_fu_369_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_375_p0 = grp_fu_369_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_375_p0 = reg_1033;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_375_p0 = grp_fu_593_p2;
        end else begin
            grp_fu_375_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_375_p1 = grp_fu_570_p2;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_375_p1 = grp_fu_589_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_375_p1 = grp_fu_603_p2;
        end else begin
            grp_fu_375_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_379_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_379_opcode = 2'd0;
        end else begin
            grp_fu_379_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_379_p0 = reg_1068;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_379_p0 = grp_fu_599_p2;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_379_p0 = grp_fu_375_p2;
        end else begin
            grp_fu_379_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_379_p1 = grp_fu_576_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_379_p1 = grp_fu_609_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_379_p1 = grp_fu_599_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_379_p1 = grp_fu_614_p2;
        end else begin
            grp_fu_379_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_384_p0 = grp_fu_379_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_384_p0 = grp_fu_624_p2;
        end else begin
            grp_fu_384_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_384_p1 = grp_fu_580_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_384_p1 = grp_fu_620_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_384_p1 = grp_fu_603_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_384_p1 = grp_fu_630_p2;
        end else begin
            grp_fu_384_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_388_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_388_opcode = 2'd0;
        end else begin
            grp_fu_388_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_388_p0 = sub23_reg_1536;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_388_p0 = reg_1039;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_388_p0 = grp_fu_384_p2;
        end else begin
            grp_fu_388_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_388_p1 = grp_fu_589_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_388_p1 = grp_fu_630_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_388_p1 = grp_fu_609_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_388_p1 = grp_fu_641_p2;
        end else begin
            grp_fu_388_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10))) begin
            grp_fu_393_p0 = grp_fu_388_p2;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_393_p0 = grp_fu_651_p2;
        end else begin
            grp_fu_393_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_393_p1 = grp_fu_593_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_393_p1 = grp_fu_657_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_393_p1 = grp_fu_614_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_393_p1 = grp_fu_661_p2;
        end else begin
            grp_fu_393_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_397_p0 = add25_reg_1541;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_397_p0 = grp_fu_624_p2;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_397_p0 = grp_fu_393_p2;
        end else begin
            grp_fu_397_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_397_p1 = grp_fu_599_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_397_p1 = grp_fu_636_p2;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_397_p1 = grp_fu_667_p2;
        end else begin
            grp_fu_397_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_402_p0 = grp_fu_651_p2;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_402_p0 = grp_fu_397_p2;
        end else begin
            grp_fu_402_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_402_p1 = grp_fu_603_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_402_p1 = grp_fu_661_p2;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_402_p1 = grp_fu_673_p2;
        end else begin
            grp_fu_402_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_411_p0 = sub28_reg_1546;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_411_p0 = grp_fu_711_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_411_p0 = grp_fu_402_p2;
        end else begin
            grp_fu_411_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_411_p1 = grp_fu_609_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_411_p1 = grp_fu_717_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_411_p1 = grp_fu_673_p2;
        end else begin
            grp_fu_411_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_416_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10))) begin
            grp_fu_416_opcode = 2'd0;
        end else begin
            grp_fu_416_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_416_p0 = grp_fu_411_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_416_p0 = grp_fu_705_p2;
        end else begin
            grp_fu_416_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_416_p1 = grp_fu_614_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_416_p1 = mul77_fu_751_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_416_p1 = grp_fu_711_p2;
        end else begin
            grp_fu_416_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_420_p0 = add33_reg_1556;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_420_p0 = grp_fu_416_p2;
        end else begin
            grp_fu_420_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_420_p1 = grp_fu_620_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_420_p1 = mul78_fu_757_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_420_p1 = grp_fu_717_p2;
        end else begin
            grp_fu_420_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_428_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_428_opcode = 2'd0;
        end else begin
            grp_fu_428_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_428_p0 = grp_fu_420_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_428_p0 = sub21_reg_1492;
        end else begin
            grp_fu_428_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_428_p1 = grp_fu_624_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_428_p1 = mul88_fu_768_p2;
        end else begin
            grp_fu_428_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_432_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_432_opcode = 2'd0;
        end else begin
            grp_fu_432_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_432_p0 = sub35_reg_1561;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_432_p0 = grp_fu_428_p2;
        end else begin
            grp_fu_432_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_432_p1 = grp_fu_630_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_432_p1 = mul89_fu_774_p2;
        end else begin
            grp_fu_432_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_437_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_437_opcode = 2'd0;
        end else begin
            grp_fu_437_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_437_p1 = grp_fu_636_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_437_p1 = mul90_fu_780_p2;
        end else begin
            grp_fu_437_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_442_p0 = add38_reg_1566;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_442_p0 = mul92_fu_790_p2;
        end else begin
            grp_fu_442_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_442_p1 = grp_fu_641_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_442_p1 = mul94_fu_801_p2;
        end else begin
            grp_fu_442_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_446_opcode = 2'd1;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_446_opcode = 2'd0;
        end else begin
            grp_fu_446_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_446_p1 = grp_fu_647_p2;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_446_p1 = mul96_fu_811_p2;
        end else begin
            grp_fu_446_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_556_p0 = mul61_reg_1509;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_556_p0 = reg_1058;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_556_p0 = m_load_10_reg_1432;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_556_p0 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_556_p0 = m_load_reg_1200;
        end else begin
            grp_fu_556_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_556_p1 = m_load_3_reg_1265;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_556_p1 = m_load_2_reg_1245;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_556_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_556_p1 = m_load_1_reg_1215;
        end else begin
            grp_fu_556_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_560_p0 = reg_1058;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_560_p0 = m_load_5_reg_1313;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_560_p0 = grp_fu_556_p2;
        end else begin
            grp_fu_560_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_560_p1 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_560_p1 = m_q1;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_560_p1 = m_load_4_reg_1292;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_560_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_560_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_566_p0 = mul71_reg_1523;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_566_p0 = grp_fu_560_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_566_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_566_p0 = m_load_8_reg_1387;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_566_p0 = m_load_reg_1200;
        end else begin
            grp_fu_566_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_566_p1 = m_load_4_reg_1292;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_566_p1 = m_load_6_reg_1342;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_566_p1 = m_load_3_reg_1265;
        end else begin
            grp_fu_566_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_570_p0 = reg_1058;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_570_p0 = m_load_8_reg_1387;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_570_p0 = grp_fu_566_p2;
        end else begin
            grp_fu_570_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_570_p1 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_570_p1 = m_load_13_reg_1483;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_570_p1 = m_load_3_reg_1265;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_570_p1 = m_load_4_reg_1292;
        end else begin
            grp_fu_570_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_576_p0 = mul71_reg_1523;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_576_p0 = grp_fu_570_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_576_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_576_p0 = m_load_8_reg_1387;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_576_p0 = m_load_5_reg_1313;
        end else begin
            grp_fu_576_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_576_p1 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_576_p1 = m_load_3_reg_1265;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_576_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_576_p1 = m_load_6_reg_1342;
        end else begin
            grp_fu_576_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_580_p0 = mul61_reg_1509;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_580_p0 = m_load_8_reg_1387;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_580_p0 = grp_fu_576_p2;
        end else begin
            grp_fu_580_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_580_p1 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_580_p1 = m_q1;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_580_p1 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_580_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_580_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_589_p0 = mul61_reg_1509;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_589_p0 = grp_fu_580_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_589_p0 = grp_fu_556_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_589_p0 = m_load_1_reg_1215;
        end else begin
            grp_fu_589_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_589_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_589_p1 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_589_p1 = m_load_8_reg_1387;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_589_p1 = bitcast_ln42_1_fu_1083_p1;
        end else begin
            grp_fu_589_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_593_p0 = reg_1058;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_593_p0 = m_q0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_593_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_593_p0 = grp_fu_589_p2;
        end else begin
            grp_fu_593_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_593_p1 = m_load_6_reg_1342;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_593_p1 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_593_p1 = m_load_reg_1200;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_593_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_593_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_599_p0 = mul71_reg_1523;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_599_p0 = grp_fu_593_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_599_p0 = m_load_9_reg_1406;
        end else begin
            grp_fu_599_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_599_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_599_p1 = m_load_2_reg_1245;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_599_p1 = m_load_3_reg_1265;
        end else begin
            grp_fu_599_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_603_p0 = reg_1058;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_603_p0 = m_q0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_603_p0 = grp_fu_576_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_603_p0 = grp_fu_599_p2;
        end else begin
            grp_fu_603_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_603_p1 = m_load_reg_1200;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_603_p1 = m_load_3_reg_1265;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_603_p1 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_603_p1 = m_load_4_reg_1292;
        end else begin
            grp_fu_603_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_609_p0 = mul71_reg_1523;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_609_p0 = grp_fu_603_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_609_p0 = grp_fu_593_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_609_p0 = m_q1;
        end else begin
            grp_fu_609_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_609_p1 = m_load_4_reg_1292;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_609_p1 = m_load_1_reg_1215;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_609_p1 = m_load_6_reg_1342;
        end else begin
            grp_fu_609_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_614_p0 = mul61_reg_1509;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_614_p0 = m_load_10_reg_1432;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_614_p0 = grp_fu_566_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_614_p0 = grp_fu_609_p2;
        end else begin
            grp_fu_614_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_614_p1 = m_load_reg_1200;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_614_p1 = m_load_13_reg_1483;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_614_p1 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_614_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_614_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_620_p0 = mul57_reg_1497;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_620_p0 = grp_fu_614_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_620_p0 = m_load_1_reg_1215;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_620_p0 = m_load_9_reg_1406;
        end else begin
            grp_fu_620_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_620_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_620_p1 = m_load_2_reg_1245;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_620_p1 = bitcast_ln63_1_fu_1099_p1;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_620_p1 = m_load_5_reg_1313;
        end else begin
            grp_fu_620_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_624_p0 = mul59_reg_1503;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_624_p0 = m_load_10_reg_1432;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_624_p0 = grp_fu_620_p2;
        end else begin
            grp_fu_624_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_624_p1 = m_load_6_reg_1342;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_624_p1 = m_q1;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_624_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_624_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_630_p0 = mul68_reg_1517;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_630_p0 = grp_fu_624_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_630_p0 = m_q1;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_630_p0 = grp_fu_599_p2;
        end else begin
            grp_fu_630_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_630_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_630_p1 = m_load_4_reg_1292;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_630_p1 = m_load_3_reg_1265;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_630_p1 = m_load_8_reg_1387;
        end else begin
            grp_fu_630_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_636_p0 = mul59_reg_1503;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_636_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_636_p0 = grp_fu_630_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_636_p0 = m_q1;
        end else begin
            grp_fu_636_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_636_p1 = m_load_13_reg_1483;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_636_p1 = m_load_4_reg_1292;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_636_p1 = m_load_reg_1200;
        end else begin
            grp_fu_636_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_641_p0 = mul68_reg_1517;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_641_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_641_p0 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_641_p0 = grp_fu_636_p2;
        end else begin
            grp_fu_641_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_641_p1 = m_load_6_reg_1342;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_641_p1 = m_q1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_641_p1 = m_q0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_641_p1 = m_load_2_reg_1245;
        end else begin
            grp_fu_641_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_647_p0 = mul57_reg_1497;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_647_p0 = m_q1;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_647_p0 = m_load_5_reg_1313;
        end else begin
            grp_fu_647_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_647_p1 = m_load_reg_1200;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_647_p1 = bitcast_ln77_1_fu_1115_p1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_647_p1 = m_load_6_reg_1342;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_647_p1 = bitcast_ln42_1_fu_1083_p1;
        end else begin
            grp_fu_647_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state9))) begin
            grp_fu_651_p1 = m_load_2_reg_1245;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_651_p1 = m_load_4_reg_1292;
        end else begin
            grp_fu_651_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_657_p0 = grp_fu_603_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_657_p0 = m_q1;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_657_p0 = m_load_9_reg_1406;
        end else begin
            grp_fu_657_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_657_p1 = m_load_8_reg_1387;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_657_p1 = m_load_7_reg_1358;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_657_p1 = m_load_1_reg_1215;
        end else begin
            grp_fu_657_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_661_p0 = m_load_10_reg_1432;
        end else if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_661_p0 = grp_fu_657_p2;
        end else begin
            grp_fu_661_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_661_p1 = m_load_12_reg_1470;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_661_p1 = m_load_4_reg_1292;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_661_p1 = m_load_8_reg_1387;
        end else begin
            grp_fu_661_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_667_p0 = grp_fu_661_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_667_p0 = m_load_reg_1200;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_667_p0 = grp_fu_636_p2;
        end else begin
            grp_fu_667_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_667_p1 = m_load_2_reg_1245;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_667_p1 = m_q0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_667_p1 = m_load_4_reg_1292;
        end else begin
            grp_fu_667_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_673_p0 = grp_fu_624_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_673_p0 = grp_fu_667_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_673_p0 = grp_fu_609_p2;
        end else begin
            grp_fu_673_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_673_p1 = m_load_2_reg_1245;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7))) begin
            grp_fu_673_p1 = m_load_8_reg_1387;
        end else begin
            grp_fu_673_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_701_p0 = m_load_11_reg_1445;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_701_p0 = m_load_6_reg_1342;
        end else begin
            grp_fu_701_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_701_p1 = m_load_12_reg_1470;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_701_p1 = bitcast_ln63_1_fu_1099_p1;
        end else begin
            grp_fu_701_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_705_p0 = m_q0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_705_p0 = grp_fu_701_p2;
        end else begin
            grp_fu_705_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_705_p1 = m_load_5_reg_1313;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_705_p1 = m_load_3_reg_1265;
        end else begin
            grp_fu_705_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_711_p0 = grp_fu_705_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_711_p0 = grp_fu_657_p2;
        end else begin
            grp_fu_711_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_711_p1 = m_load_4_reg_1292;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_711_p1 = m_load_1_reg_1215;
        end else begin
            grp_fu_711_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_717_p0 = grp_fu_593_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_717_p0 = grp_fu_667_p2;
        end else begin
            grp_fu_717_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_717_p1 = m_load_8_reg_1387;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_717_p1 = m_load_3_reg_1265;
        end else begin
            grp_fu_717_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state14)) begin
            inv_address0 = 64'd7;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            inv_address0 = 64'd14;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            inv_address0 = 64'd6;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            inv_address0 = 64'd13;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            inv_address0 = 64'd5;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            inv_address0 = 64'd12;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            inv_address0 = 64'd8;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            inv_address0 = 64'd0;
        end else if (((1'd0 == and_ln149_reg_1597) & (1'b1 == ap_CS_fsm_state17))) begin
            inv_address0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_address0;
        end else begin
            inv_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            inv_address1 = 64'd15;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            inv_address1 = 64'd11;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            inv_address1 = 64'd3;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            inv_address1 = 64'd10;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            inv_address1 = 64'd2;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            inv_address1 = 64'd9;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            inv_address1 = 64'd1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            inv_address1 = 64'd4;
        end else begin
            inv_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11))) begin
            inv_ce0 = 1'b1;
        end else if (((1'd0 == and_ln149_reg_1597) & (1'b1 == ap_CS_fsm_state17))) begin
            inv_ce0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_inv_ce0;
        end else begin
            inv_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state15))) begin
            inv_ce1 = 1'b1;
        end else begin
            inv_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state14)) begin
            inv_d0 = sub34_reg_1582;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            inv_d0 = add29_reg_1577;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            inv_d0 = reg_1046;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            inv_d0 = grp_fu_364_p2;
        end else if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state12))) begin
            inv_d0 = reg_1052;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            inv_d0 = grp_fu_384_p2;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            inv_d0 = grp_fu_369_p2;
        end else begin
            inv_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            inv_d1 = sub39_reg_1592;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            inv_d1 = add37_reg_1587;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            inv_d1 = add32_reg_1551;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            inv_d1 = reg_1039;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            inv_d1 = sub22_reg_1531;
        end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
            inv_d1 = grp_fu_375_p2;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            inv_d1 = grp_fu_369_p2;
        end else begin
            inv_d1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11))) begin
            inv_we0 = 1'b1;
        end else begin
            inv_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state15))) begin
            inv_we1 = 1'b1;
        end else begin
            inv_we1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            m_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            m_address0 = 64'd2;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            m_address0 = 64'd12;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            m_address0 = 64'd4;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            m_address0 = 64'd7;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            m_address0 = 64'd9;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            m_address0 = 64'd11;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            m_address0 = 64'd10;
        end else begin
            m_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            m_address1 = 64'd3;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            m_address1 = 64'd1;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            m_address1 = 64'd8;
        end else if ((1'b1 == ap_CS_fsm_state5)) begin
            m_address1 = 64'd13;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            m_address1 = 64'd6;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            m_address1 = 64'd14;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            m_address1 = 64'd15;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            m_address1 = 64'd5;
        end else begin
            m_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
            m_ce0 = 1'b1;
        end else begin
            m_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
            m_ce1 = 1'b1;
        end else begin
            m_ce1 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                if (((1'd1 == and_ln149_fu_1174_p2) & (1'b1 == ap_CS_fsm_state15))) begin
                    ap_NS_fsm = ap_ST_fsm_state17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state16;
                end
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                if (((1'b0 == ap_block_state17_on_subcall_done) & (1'b1 == ap_CS_fsm_state17))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state17;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign and_ln149_fu_1174_p2 = (tmp_3_fu_1028_p2 & or_ln149_fu_1168_p2);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    always @(*) begin
        ap_block_state17_on_subcall_done = ((1'd0 == and_ln149_reg_1597) & (grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_done == 1'b0));
    end

    assign bitcast_ln42_1_fu_1083_p1 = xor_ln42_fu_1077_p2;

    assign bitcast_ln42_fu_1074_p1 = m_load_9_reg_1406;

    assign bitcast_ln63_1_fu_1099_p1 = xor_ln63_fu_1093_p2;

    assign bitcast_ln63_fu_1089_p1 = m_q1;

    assign bitcast_ln77_1_fu_1115_p1 = xor_ln77_fu_1109_p2;

    assign bitcast_ln77_fu_1105_p1 = m_q0;

    assign data_fu_1122_p1 = det_2_reg_1571;

    assign grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_ap_start_reg;

    assign icmp_ln149_1_fu_1162_p2 = ((trunc_ln149_fu_1129_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln149_fu_1156_p2 = ((tmp_2_fu_1146_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign invOut_address0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_address0;

    assign invOut_ce0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_ce0;

    assign invOut_d0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_d0;

    assign invOut_we0 = grp_invert4x4Matrix_double_Pipeline_VITIS_LOOP_153_1_VITIS_LOOP_154_2_fu_352_invOut_we0;

    assign or_ln149_fu_1168_p2 = (icmp_ln149_fu_1156_p2 | icmp_ln149_1_fu_1162_p2);

    assign t_fu_1133_p3 = {{1'd0}, {trunc_ln479_fu_1125_p1}};

    assign tmp_2_fu_1146_p4 = {{data_fu_1122_p1[62:52]}};

    assign tmp_3_fu_1028_p0 = t_fu_1133_p3;

    assign trunc_ln149_fu_1129_p1 = data_fu_1122_p1[51:0];

    assign trunc_ln479_fu_1125_p1 = data_fu_1122_p1[62:0];

    assign xor_ln42_fu_1077_p2 = (bitcast_ln42_fu_1074_p1 ^ 64'd9223372036854775808);

    assign xor_ln63_fu_1093_p2 = (bitcast_ln63_fu_1089_p1 ^ 64'd9223372036854775808);

    assign xor_ln77_fu_1109_p2 = (bitcast_ln77_fu_1105_p1 ^ 64'd9223372036854775808);

endmodule  //main_invert4x4Matrix_double_s
