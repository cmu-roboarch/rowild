/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module main_pf_RAM_AUTO_1R1W (

    address0,
    ce0,
    d0,
    we0,
    q0,

    address1,
    ce1,
    d1,
    we1,
    q1,

    reset,
    clk
);

    parameter DataWidth = 256;
    parameter AddressWidth = 17;
    parameter AddressRange = 80504;
    parameter COL_WIDTH = 8;
    parameter NUM_COL = (DataWidth / COL_WIDTH);

    input [AddressWidth-1:0] address0;
    input ce0;
    input [DataWidth-1:0] d0;
    input [NUM_COL-1:0] we0;
    output reg [DataWidth-1:0] q0;

    input [AddressWidth-1:0] address1;
    input ce1;
    input [DataWidth-1:0] d1;
    input [NUM_COL-1:0] we1;
    output reg [DataWidth-1:0] q1;

    input reset;
    input clk;

    (* ram_style = "auto"  *) reg [DataWidth-1:0] ram[0:AddressRange-1];


    genvar i;







    //read first
    generate
        for (i = 0; i < NUM_COL; i = i + 1) begin
            always @(posedge clk) begin
                if (ce0) begin
                    if (we0[i]) begin
                        ram[address0][i*COL_WIDTH+:COL_WIDTH] <= d0[i*COL_WIDTH+:COL_WIDTH];
                    end
                    q0[i*COL_WIDTH+:COL_WIDTH] <= ram[address0][i*COL_WIDTH+:COL_WIDTH];
                end
            end
        end
    endgenerate







    //read first
    generate
        for (i = 0; i < NUM_COL; i = i + 1) begin
            always @(posedge clk) begin
                if (ce1) begin
                    if (we1[i]) begin
                        ram[address1][i*COL_WIDTH+:COL_WIDTH] <= d1[i*COL_WIDTH+:COL_WIDTH];
                    end
                    q1[i*COL_WIDTH+:COL_WIDTH] <= ram[address1][i*COL_WIDTH+:COL_WIDTH];
                end
            end
        end
    endgenerate



endmodule

