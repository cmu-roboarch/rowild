/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_2 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    empty,
    l_cPoints_address0,
    l_cPoints_ce0,
    l_cPoints_we0,
    l_cPoints_d0
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [4:0] empty;
    output [6:0] l_cPoints_address0;
    output l_cPoints_ce0;
    output l_cPoints_we0;
    output [63:0] l_cPoints_d0;

    reg ap_idle;
    reg l_cPoints_ce0;
    reg l_cPoints_we0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] exitcond238_fu_100_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire   [6:0] empty_78_fu_190_p2;
    reg   [6:0] empty_78_reg_239;
    wire    ap_block_pp0_stage0_11001;
    wire   [63:0] p_cast_fu_211_p1;
    wire    ap_block_pp0_stage0;
    reg   [4:0] phi_urem_fu_46;
    wire   [4:0] idx_urem_fu_130_p3;
    wire    ap_loop_init;
    reg   [4:0] ap_sig_allocacmp_phi_urem_load;
    reg   [10:0] phi_mul_fu_50;
    wire   [10:0] next_mul_fu_138_p2;
    reg   [10:0] ap_sig_allocacmp_phi_mul_load;
    reg   [4:0] empty_72_fu_54;
    wire   [4:0] empty_73_fu_106_p2;
    reg   [4:0] ap_sig_allocacmp_p_load;
    wire   [4:0] next_urem_fu_118_p2;
    wire   [0:0] empty_74_fu_124_p2;
    wire   [3:0] tmp_22_fu_144_p4;
    wire   [5:0] p_cast1_fu_78_p1;
    wire   [5:0] tmp_39_cast_fu_154_p1;
    wire   [5:0] empty_75_fu_158_p2;
    wire   [4:0] empty_76_fu_168_p1;
    wire   [6:0] tmp_23_fu_172_p3;
    wire   [6:0] p_cast2_fu_164_p1;
    wire   [6:0] empty_77_fu_180_p2;
    wire   [6:0] phi_urem_cast_fu_186_p1;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 phi_urem_fu_46 = 5'd0;
        #0 phi_mul_fu_50 = 11'd0;
        #0 empty_72_fu_54 = 5'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((exitcond238_fu_100_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                empty_72_fu_54 <= empty_73_fu_106_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                empty_72_fu_54 <= 5'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((exitcond238_fu_100_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                phi_mul_fu_50 <= next_mul_fu_138_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                phi_mul_fu_50 <= 11'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((exitcond238_fu_100_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                phi_urem_fu_46 <= idx_urem_fu_130_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                phi_urem_fu_46 <= 5'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            empty_78_reg_239 <= empty_78_fu_190_p2;
        end
    end

    always @(*) begin
        if (((exitcond238_fu_100_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_p_load = 5'd0;
        end else begin
            ap_sig_allocacmp_p_load = empty_72_fu_54;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_phi_mul_load = 11'd0;
        end else begin
            ap_sig_allocacmp_phi_mul_load = phi_mul_fu_50;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_phi_urem_load = 5'd0;
        end else begin
            ap_sig_allocacmp_phi_urem_load = phi_urem_fu_46;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_cPoints_ce0 = 1'b1;
        end else begin
            l_cPoints_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_cPoints_we0 = 1'b1;
        end else begin
            l_cPoints_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign empty_73_fu_106_p2 = (ap_sig_allocacmp_p_load + 5'd1);

    assign empty_74_fu_124_p2 = ((next_urem_fu_118_p2 < 5'd3) ? 1'b1 : 1'b0);

    assign empty_75_fu_158_p2 = (p_cast1_fu_78_p1 + tmp_39_cast_fu_154_p1);

    assign empty_76_fu_168_p1 = empty_75_fu_158_p2[4:0];

    assign empty_77_fu_180_p2 = (tmp_23_fu_172_p3 - p_cast2_fu_164_p1);

    assign empty_78_fu_190_p2 = (empty_77_fu_180_p2 + phi_urem_cast_fu_186_p1);

    assign exitcond238_fu_100_p2 = ((ap_sig_allocacmp_p_load == 5'd27) ? 1'b1 : 1'b0);

    assign idx_urem_fu_130_p3 = ((empty_74_fu_124_p2[0:0] == 1'b1) ? next_urem_fu_118_p2 : 5'd0);

    assign l_cPoints_address0 = p_cast_fu_211_p1;

    assign l_cPoints_d0 = 64'd0;

    assign next_mul_fu_138_p2 = (ap_sig_allocacmp_phi_mul_load + 11'd43);

    assign next_urem_fu_118_p2 = (ap_sig_allocacmp_phi_urem_load + 5'd1);

    assign p_cast1_fu_78_p1 = empty;

    assign p_cast2_fu_164_p1 = empty_75_fu_158_p2;

    assign p_cast_fu_211_p1 = empty_78_reg_239;

    assign phi_urem_cast_fu_186_p1 = ap_sig_allocacmp_phi_urem_load;

    assign tmp_22_fu_144_p4 = {{ap_sig_allocacmp_phi_mul_load[10:7]}};

    assign tmp_23_fu_172_p3 = {{empty_76_fu_168_p1}, {2'd0}};

    assign tmp_39_cast_fu_154_p1 = tmp_22_fu_144_p4;

endmodule  //main_main_Pipeline_2
