/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_updateMotion (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    pf_address0,
    pf_ce0,
    pf_we0,
    pf_d0,
    pf_q0,
    prevOdometry_0_0_val,
    prevOdometry_0_1_val,
    prevOdometry_0_2_val,
    currOdometry_0_0_val,
    currOdometry_0_1_val,
    currOdometry_0_2_val,
    grp_fu_394_p_din0,
    grp_fu_394_p_dout0,
    grp_fu_394_p_ce,
    grp_fu_397_p_din0,
    grp_fu_397_p_din1,
    grp_fu_397_p_opcode,
    grp_fu_397_p_dout0,
    grp_fu_397_p_ce,
    grp_fu_401_p_din0,
    grp_fu_401_p_din1,
    grp_fu_401_p_opcode,
    grp_fu_401_p_dout0,
    grp_fu_401_p_ce,
    grp_fu_405_p_din0,
    grp_fu_405_p_din1,
    grp_fu_405_p_dout0,
    grp_fu_405_p_ce,
    grp_fu_409_p_din0,
    grp_fu_409_p_din1,
    grp_fu_409_p_dout0,
    grp_fu_409_p_ce,
    grp_fu_413_p_din0,
    grp_fu_413_p_din1,
    grp_fu_413_p_opcode,
    grp_fu_413_p_dout0,
    grp_fu_413_p_ce,
    grp_fu_417_p_din0,
    grp_fu_417_p_din1,
    grp_fu_417_p_dout0,
    grp_fu_417_p_ce,
    grp_sin_or_cos_double_s_fu_421_p_din1,
    grp_sin_or_cos_double_s_fu_421_p_din2,
    grp_sin_or_cos_double_s_fu_421_p_dout0,
    grp_sin_or_cos_double_s_fu_421_p_start,
    grp_sin_or_cos_double_s_fu_421_p_ready,
    grp_sin_or_cos_double_s_fu_421_p_done,
    grp_sin_or_cos_double_s_fu_421_p_idle,
    grp_sin_or_cos_double_s_fu_432_p_din1,
    grp_sin_or_cos_double_s_fu_432_p_din2,
    grp_sin_or_cos_double_s_fu_432_p_dout0,
    grp_sin_or_cos_double_s_fu_432_p_start,
    grp_sin_or_cos_double_s_fu_432_p_ready,
    grp_sin_or_cos_double_s_fu_432_p_done,
    grp_sin_or_cos_double_s_fu_432_p_idle
);

    parameter ap_ST_fsm_state1 = 243'd1;
    parameter ap_ST_fsm_state2 = 243'd2;
    parameter ap_ST_fsm_state3 = 243'd4;
    parameter ap_ST_fsm_state4 = 243'd8;
    parameter ap_ST_fsm_state5 = 243'd16;
    parameter ap_ST_fsm_state6 = 243'd32;
    parameter ap_ST_fsm_state7 = 243'd64;
    parameter ap_ST_fsm_state8 = 243'd128;
    parameter ap_ST_fsm_state9 = 243'd256;
    parameter ap_ST_fsm_state10 = 243'd512;
    parameter ap_ST_fsm_state11 = 243'd1024;
    parameter ap_ST_fsm_state12 = 243'd2048;
    parameter ap_ST_fsm_state13 = 243'd4096;
    parameter ap_ST_fsm_state14 = 243'd8192;
    parameter ap_ST_fsm_state15 = 243'd16384;
    parameter ap_ST_fsm_state16 = 243'd32768;
    parameter ap_ST_fsm_state17 = 243'd65536;
    parameter ap_ST_fsm_state18 = 243'd131072;
    parameter ap_ST_fsm_state19 = 243'd262144;
    parameter ap_ST_fsm_state20 = 243'd524288;
    parameter ap_ST_fsm_state21 = 243'd1048576;
    parameter ap_ST_fsm_state22 = 243'd2097152;
    parameter ap_ST_fsm_state23 = 243'd4194304;
    parameter ap_ST_fsm_state24 = 243'd8388608;
    parameter ap_ST_fsm_state25 = 243'd16777216;
    parameter ap_ST_fsm_state26 = 243'd33554432;
    parameter ap_ST_fsm_state27 = 243'd67108864;
    parameter ap_ST_fsm_state28 = 243'd134217728;
    parameter ap_ST_fsm_state29 = 243'd268435456;
    parameter ap_ST_fsm_state30 = 243'd536870912;
    parameter ap_ST_fsm_state31 = 243'd1073741824;
    parameter ap_ST_fsm_state32 = 243'd2147483648;
    parameter ap_ST_fsm_state33 = 243'd4294967296;
    parameter ap_ST_fsm_state34 = 243'd8589934592;
    parameter ap_ST_fsm_state35 = 243'd17179869184;
    parameter ap_ST_fsm_state36 = 243'd34359738368;
    parameter ap_ST_fsm_state37 = 243'd68719476736;
    parameter ap_ST_fsm_state38 = 243'd137438953472;
    parameter ap_ST_fsm_state39 = 243'd274877906944;
    parameter ap_ST_fsm_state40 = 243'd549755813888;
    parameter ap_ST_fsm_state41 = 243'd1099511627776;
    parameter ap_ST_fsm_state42 = 243'd2199023255552;
    parameter ap_ST_fsm_state43 = 243'd4398046511104;
    parameter ap_ST_fsm_state44 = 243'd8796093022208;
    parameter ap_ST_fsm_state45 = 243'd17592186044416;
    parameter ap_ST_fsm_state46 = 243'd35184372088832;
    parameter ap_ST_fsm_state47 = 243'd70368744177664;
    parameter ap_ST_fsm_state48 = 243'd140737488355328;
    parameter ap_ST_fsm_state49 = 243'd281474976710656;
    parameter ap_ST_fsm_state50 = 243'd562949953421312;
    parameter ap_ST_fsm_state51 = 243'd1125899906842624;
    parameter ap_ST_fsm_state52 = 243'd2251799813685248;
    parameter ap_ST_fsm_state53 = 243'd4503599627370496;
    parameter ap_ST_fsm_state54 = 243'd9007199254740992;
    parameter ap_ST_fsm_state55 = 243'd18014398509481984;
    parameter ap_ST_fsm_state56 = 243'd36028797018963968;
    parameter ap_ST_fsm_state57 = 243'd72057594037927936;
    parameter ap_ST_fsm_state58 = 243'd144115188075855872;
    parameter ap_ST_fsm_state59 = 243'd288230376151711744;
    parameter ap_ST_fsm_state60 = 243'd576460752303423488;
    parameter ap_ST_fsm_state61 = 243'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 243'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 243'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 243'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 243'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 243'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 243'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 243'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 243'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 243'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 243'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 243'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 243'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 243'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 243'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 243'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 243'd75557863725914323419136;
    parameter ap_ST_fsm_state78 = 243'd151115727451828646838272;
    parameter ap_ST_fsm_state79 = 243'd302231454903657293676544;
    parameter ap_ST_fsm_state80 = 243'd604462909807314587353088;
    parameter ap_ST_fsm_state81 = 243'd1208925819614629174706176;
    parameter ap_ST_fsm_state82 = 243'd2417851639229258349412352;
    parameter ap_ST_fsm_state83 = 243'd4835703278458516698824704;
    parameter ap_ST_fsm_state84 = 243'd9671406556917033397649408;
    parameter ap_ST_fsm_state85 = 243'd19342813113834066795298816;
    parameter ap_ST_fsm_state86 = 243'd38685626227668133590597632;
    parameter ap_ST_fsm_state87 = 243'd77371252455336267181195264;
    parameter ap_ST_fsm_state88 = 243'd154742504910672534362390528;
    parameter ap_ST_fsm_state89 = 243'd309485009821345068724781056;
    parameter ap_ST_fsm_state90 = 243'd618970019642690137449562112;
    parameter ap_ST_fsm_state91 = 243'd1237940039285380274899124224;
    parameter ap_ST_fsm_state92 = 243'd2475880078570760549798248448;
    parameter ap_ST_fsm_state93 = 243'd4951760157141521099596496896;
    parameter ap_ST_fsm_state94 = 243'd9903520314283042199192993792;
    parameter ap_ST_fsm_state95 = 243'd19807040628566084398385987584;
    parameter ap_ST_fsm_state96 = 243'd39614081257132168796771975168;
    parameter ap_ST_fsm_state97 = 243'd79228162514264337593543950336;
    parameter ap_ST_fsm_state98 = 243'd158456325028528675187087900672;
    parameter ap_ST_fsm_state99 = 243'd316912650057057350374175801344;
    parameter ap_ST_fsm_state100 = 243'd633825300114114700748351602688;
    parameter ap_ST_fsm_state101 = 243'd1267650600228229401496703205376;
    parameter ap_ST_fsm_state102 = 243'd2535301200456458802993406410752;
    parameter ap_ST_fsm_state103 = 243'd5070602400912917605986812821504;
    parameter ap_ST_fsm_state104 = 243'd10141204801825835211973625643008;
    parameter ap_ST_fsm_state105 = 243'd20282409603651670423947251286016;
    parameter ap_ST_fsm_state106 = 243'd40564819207303340847894502572032;
    parameter ap_ST_fsm_state107 = 243'd81129638414606681695789005144064;
    parameter ap_ST_fsm_state108 = 243'd162259276829213363391578010288128;
    parameter ap_ST_fsm_state109 = 243'd324518553658426726783156020576256;
    parameter ap_ST_fsm_state110 = 243'd649037107316853453566312041152512;
    parameter ap_ST_fsm_state111 = 243'd1298074214633706907132624082305024;
    parameter ap_ST_fsm_state112 = 243'd2596148429267413814265248164610048;
    parameter ap_ST_fsm_state113 = 243'd5192296858534827628530496329220096;
    parameter ap_ST_fsm_state114 = 243'd10384593717069655257060992658440192;
    parameter ap_ST_fsm_state115 = 243'd20769187434139310514121985316880384;
    parameter ap_ST_fsm_state116 = 243'd41538374868278621028243970633760768;
    parameter ap_ST_fsm_state117 = 243'd83076749736557242056487941267521536;
    parameter ap_ST_fsm_state118 = 243'd166153499473114484112975882535043072;
    parameter ap_ST_fsm_state119 = 243'd332306998946228968225951765070086144;
    parameter ap_ST_fsm_state120 = 243'd664613997892457936451903530140172288;
    parameter ap_ST_fsm_state121 = 243'd1329227995784915872903807060280344576;
    parameter ap_ST_fsm_state122 = 243'd2658455991569831745807614120560689152;
    parameter ap_ST_fsm_state123 = 243'd5316911983139663491615228241121378304;
    parameter ap_ST_fsm_state124 = 243'd10633823966279326983230456482242756608;
    parameter ap_ST_fsm_state125 = 243'd21267647932558653966460912964485513216;
    parameter ap_ST_fsm_state126 = 243'd42535295865117307932921825928971026432;
    parameter ap_ST_fsm_state127 = 243'd85070591730234615865843651857942052864;
    parameter ap_ST_fsm_state128 = 243'd170141183460469231731687303715884105728;
    parameter ap_ST_fsm_state129 = 243'd340282366920938463463374607431768211456;
    parameter ap_ST_fsm_state130 = 243'd680564733841876926926749214863536422912;
    parameter ap_ST_fsm_state131 = 243'd1361129467683753853853498429727072845824;
    parameter ap_ST_fsm_state132 = 243'd2722258935367507707706996859454145691648;
    parameter ap_ST_fsm_state133 = 243'd5444517870735015415413993718908291383296;
    parameter ap_ST_fsm_state134 = 243'd10889035741470030830827987437816582766592;
    parameter ap_ST_fsm_state135 = 243'd21778071482940061661655974875633165533184;
    parameter ap_ST_fsm_state136 = 243'd43556142965880123323311949751266331066368;
    parameter ap_ST_fsm_state137 = 243'd87112285931760246646623899502532662132736;
    parameter ap_ST_fsm_state138 = 243'd174224571863520493293247799005065324265472;
    parameter ap_ST_fsm_state139 = 243'd348449143727040986586495598010130648530944;
    parameter ap_ST_fsm_state140 = 243'd696898287454081973172991196020261297061888;
    parameter ap_ST_fsm_state141 = 243'd1393796574908163946345982392040522594123776;
    parameter ap_ST_fsm_state142 = 243'd2787593149816327892691964784081045188247552;
    parameter ap_ST_fsm_state143 = 243'd5575186299632655785383929568162090376495104;
    parameter ap_ST_fsm_state144 = 243'd11150372599265311570767859136324180752990208;
    parameter ap_ST_fsm_state145 = 243'd22300745198530623141535718272648361505980416;
    parameter ap_ST_fsm_state146 = 243'd44601490397061246283071436545296723011960832;
    parameter ap_ST_fsm_state147 = 243'd89202980794122492566142873090593446023921664;
    parameter ap_ST_fsm_state148 = 243'd178405961588244985132285746181186892047843328;
    parameter ap_ST_fsm_state149 = 243'd356811923176489970264571492362373784095686656;
    parameter ap_ST_fsm_state150 = 243'd713623846352979940529142984724747568191373312;
    parameter ap_ST_fsm_state151 = 243'd1427247692705959881058285969449495136382746624;
    parameter ap_ST_fsm_state152 = 243'd2854495385411919762116571938898990272765493248;
    parameter ap_ST_fsm_state153 = 243'd5708990770823839524233143877797980545530986496;
    parameter ap_ST_fsm_state154 = 243'd11417981541647679048466287755595961091061972992;
    parameter ap_ST_fsm_state155 = 243'd22835963083295358096932575511191922182123945984;
    parameter ap_ST_fsm_state156 = 243'd45671926166590716193865151022383844364247891968;
    parameter ap_ST_fsm_state157 = 243'd91343852333181432387730302044767688728495783936;
    parameter ap_ST_fsm_state158 = 243'd182687704666362864775460604089535377456991567872;
    parameter ap_ST_fsm_state159 = 243'd365375409332725729550921208179070754913983135744;
    parameter ap_ST_fsm_state160 = 243'd730750818665451459101842416358141509827966271488;
    parameter ap_ST_fsm_state161 = 243'd1461501637330902918203684832716283019655932542976;
    parameter ap_ST_fsm_state162 = 243'd2923003274661805836407369665432566039311865085952;
    parameter ap_ST_fsm_state163 = 243'd5846006549323611672814739330865132078623730171904;
    parameter ap_ST_fsm_state164 = 243'd11692013098647223345629478661730264157247460343808;
    parameter ap_ST_fsm_state165 = 243'd23384026197294446691258957323460528314494920687616;
    parameter ap_ST_fsm_state166 = 243'd46768052394588893382517914646921056628989841375232;
    parameter ap_ST_fsm_state167 = 243'd93536104789177786765035829293842113257979682750464;
    parameter ap_ST_fsm_state168 = 243'd187072209578355573530071658587684226515959365500928;
    parameter ap_ST_fsm_state169 = 243'd374144419156711147060143317175368453031918731001856;
    parameter ap_ST_fsm_state170 = 243'd748288838313422294120286634350736906063837462003712;
    parameter ap_ST_fsm_state171 = 243'd1496577676626844588240573268701473812127674924007424;
    parameter ap_ST_fsm_state172 = 243'd2993155353253689176481146537402947624255349848014848;
    parameter ap_ST_fsm_state173 = 243'd5986310706507378352962293074805895248510699696029696;
    parameter ap_ST_fsm_state174 = 243'd11972621413014756705924586149611790497021399392059392;
    parameter ap_ST_fsm_state175 = 243'd23945242826029513411849172299223580994042798784118784;
    parameter ap_ST_fsm_state176 = 243'd47890485652059026823698344598447161988085597568237568;
    parameter ap_ST_fsm_state177 = 243'd95780971304118053647396689196894323976171195136475136;
    parameter ap_ST_fsm_state178 = 243'd191561942608236107294793378393788647952342390272950272;
    parameter ap_ST_fsm_state179 = 243'd383123885216472214589586756787577295904684780545900544;
    parameter ap_ST_fsm_state180 = 243'd766247770432944429179173513575154591809369561091801088;
    parameter ap_ST_fsm_state181 = 243'd1532495540865888858358347027150309183618739122183602176;
    parameter ap_ST_fsm_state182 = 243'd3064991081731777716716694054300618367237478244367204352;
    parameter ap_ST_fsm_state183 = 243'd6129982163463555433433388108601236734474956488734408704;
    parameter ap_ST_fsm_state184 = 243'd12259964326927110866866776217202473468949912977468817408;
    parameter ap_ST_fsm_state185 = 243'd24519928653854221733733552434404946937899825954937634816;
    parameter ap_ST_fsm_state186 = 243'd49039857307708443467467104868809893875799651909875269632;
    parameter ap_ST_fsm_state187 = 243'd98079714615416886934934209737619787751599303819750539264;
    parameter ap_ST_fsm_state188 = 243'd196159429230833773869868419475239575503198607639501078528;
    parameter ap_ST_fsm_state189 = 243'd392318858461667547739736838950479151006397215279002157056;
    parameter ap_ST_fsm_state190 = 243'd784637716923335095479473677900958302012794430558004314112;
    parameter ap_ST_fsm_state191 = 243'd1569275433846670190958947355801916604025588861116008628224;
    parameter ap_ST_fsm_state192 = 243'd3138550867693340381917894711603833208051177722232017256448;
    parameter ap_ST_fsm_state193 = 243'd6277101735386680763835789423207666416102355444464034512896;
    parameter ap_ST_fsm_state194 = 243'd12554203470773361527671578846415332832204710888928069025792;
    parameter ap_ST_fsm_state195 = 243'd25108406941546723055343157692830665664409421777856138051584;
    parameter ap_ST_fsm_state196 = 243'd50216813883093446110686315385661331328818843555712276103168;
    parameter    ap_ST_fsm_state197 = 243'd100433627766186892221372630771322662657637687111424552206336;
    parameter    ap_ST_fsm_state198 = 243'd200867255532373784442745261542645325315275374222849104412672;
    parameter    ap_ST_fsm_state199 = 243'd401734511064747568885490523085290650630550748445698208825344;
    parameter    ap_ST_fsm_state200 = 243'd803469022129495137770981046170581301261101496891396417650688;
    parameter    ap_ST_fsm_state201 = 243'd1606938044258990275541962092341162602522202993782792835301376;
    parameter    ap_ST_fsm_state202 = 243'd3213876088517980551083924184682325205044405987565585670602752;
    parameter    ap_ST_fsm_state203 = 243'd6427752177035961102167848369364650410088811975131171341205504;
    parameter    ap_ST_fsm_state204 = 243'd12855504354071922204335696738729300820177623950262342682411008;
    parameter    ap_ST_fsm_state205 = 243'd25711008708143844408671393477458601640355247900524685364822016;
    parameter    ap_ST_fsm_state206 = 243'd51422017416287688817342786954917203280710495801049370729644032;
    parameter    ap_ST_fsm_state207 = 243'd102844034832575377634685573909834406561420991602098741459288064;
    parameter    ap_ST_fsm_state208 = 243'd205688069665150755269371147819668813122841983204197482918576128;
    parameter    ap_ST_fsm_state209 = 243'd411376139330301510538742295639337626245683966408394965837152256;
    parameter    ap_ST_fsm_state210 = 243'd822752278660603021077484591278675252491367932816789931674304512;
    parameter    ap_ST_fsm_state211 = 243'd1645504557321206042154969182557350504982735865633579863348609024;
    parameter    ap_ST_fsm_state212 = 243'd3291009114642412084309938365114701009965471731267159726697218048;
    parameter    ap_ST_fsm_state213 = 243'd6582018229284824168619876730229402019930943462534319453394436096;
    parameter    ap_ST_fsm_state214 = 243'd13164036458569648337239753460458804039861886925068638906788872192;
    parameter    ap_ST_fsm_state215 = 243'd26328072917139296674479506920917608079723773850137277813577744384;
    parameter    ap_ST_fsm_state216 = 243'd52656145834278593348959013841835216159447547700274555627155488768;
    parameter    ap_ST_fsm_state217 = 243'd105312291668557186697918027683670432318895095400549111254310977536;
    parameter    ap_ST_fsm_state218 = 243'd210624583337114373395836055367340864637790190801098222508621955072;
    parameter    ap_ST_fsm_state219 = 243'd421249166674228746791672110734681729275580381602196445017243910144;
    parameter    ap_ST_fsm_state220 = 243'd842498333348457493583344221469363458551160763204392890034487820288;
    parameter    ap_ST_fsm_state221 = 243'd1684996666696914987166688442938726917102321526408785780068975640576;
    parameter    ap_ST_fsm_state222 = 243'd3369993333393829974333376885877453834204643052817571560137951281152;
    parameter    ap_ST_fsm_state223 = 243'd6739986666787659948666753771754907668409286105635143120275902562304;
    parameter    ap_ST_fsm_state224 = 243'd13479973333575319897333507543509815336818572211270286240551805124608;
    parameter    ap_ST_fsm_state225 = 243'd26959946667150639794667015087019630673637144422540572481103610249216;
    parameter    ap_ST_fsm_state226 = 243'd53919893334301279589334030174039261347274288845081144962207220498432;
    parameter    ap_ST_fsm_state227 = 243'd107839786668602559178668060348078522694548577690162289924414440996864;
    parameter    ap_ST_fsm_state228 = 243'd215679573337205118357336120696157045389097155380324579848828881993728;
    parameter    ap_ST_fsm_state229 = 243'd431359146674410236714672241392314090778194310760649159697657763987456;
    parameter    ap_ST_fsm_state230 = 243'd862718293348820473429344482784628181556388621521298319395315527974912;
    parameter    ap_ST_fsm_state231 = 243'd1725436586697640946858688965569256363112777243042596638790631055949824;
    parameter    ap_ST_fsm_state232 = 243'd3450873173395281893717377931138512726225554486085193277581262111899648;
    parameter    ap_ST_fsm_state233 = 243'd6901746346790563787434755862277025452451108972170386555162524223799296;
    parameter    ap_ST_fsm_state234 = 243'd13803492693581127574869511724554050904902217944340773110325048447598592;
    parameter    ap_ST_fsm_state235 = 243'd27606985387162255149739023449108101809804435888681546220650096895197184;
    parameter    ap_ST_fsm_state236 = 243'd55213970774324510299478046898216203619608871777363092441300193790394368;
    parameter    ap_ST_fsm_state237 = 243'd110427941548649020598956093796432407239217743554726184882600387580788736;
    parameter    ap_ST_fsm_state238 = 243'd220855883097298041197912187592864814478435487109452369765200775161577472;
    parameter    ap_ST_fsm_state239 = 243'd441711766194596082395824375185729628956870974218904739530401550323154944;
    parameter    ap_ST_fsm_state240 = 243'd883423532389192164791648750371459257913741948437809479060803100646309888;
    parameter    ap_ST_fsm_state241 = 243'd1766847064778384329583297500742918515827483896875618958121606201292619776;
    parameter    ap_ST_fsm_state242 = 243'd3533694129556768659166595001485837031654967793751237916243212402585239552;
    parameter    ap_ST_fsm_state243 = 243'd7067388259113537318333190002971674063309935587502475832486424805170479104;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [16:0] pf_address0;
    output pf_ce0;
    output [31:0] pf_we0;
    output [255:0] pf_d0;
    input [255:0] pf_q0;
    input [31:0] prevOdometry_0_0_val;
    input [31:0] prevOdometry_0_1_val;
    input [31:0] prevOdometry_0_2_val;
    input [31:0] currOdometry_0_0_val;
    input [31:0] currOdometry_0_1_val;
    input [31:0] currOdometry_0_2_val;
    output [31:0] grp_fu_394_p_din0;
    input [63:0] grp_fu_394_p_dout0;
    output grp_fu_394_p_ce;
    output [63:0] grp_fu_397_p_din0;
    output [63:0] grp_fu_397_p_din1;
    output [1:0] grp_fu_397_p_opcode;
    input [63:0] grp_fu_397_p_dout0;
    output grp_fu_397_p_ce;
    output [63:0] grp_fu_401_p_din0;
    output [63:0] grp_fu_401_p_din1;
    output [1:0] grp_fu_401_p_opcode;
    input [63:0] grp_fu_401_p_dout0;
    output grp_fu_401_p_ce;
    output [63:0] grp_fu_405_p_din0;
    output [63:0] grp_fu_405_p_din1;
    input [63:0] grp_fu_405_p_dout0;
    output grp_fu_405_p_ce;
    output [63:0] grp_fu_409_p_din0;
    output [63:0] grp_fu_409_p_din1;
    input [63:0] grp_fu_409_p_dout0;
    output grp_fu_409_p_ce;
    output [63:0] grp_fu_413_p_din0;
    output [63:0] grp_fu_413_p_din1;
    output [4:0] grp_fu_413_p_opcode;
    input [0:0] grp_fu_413_p_dout0;
    output grp_fu_413_p_ce;
    output [63:0] grp_fu_417_p_din0;
    output [63:0] grp_fu_417_p_din1;
    input [63:0] grp_fu_417_p_dout0;
    output grp_fu_417_p_ce;
    output [63:0] grp_sin_or_cos_double_s_fu_421_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_421_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_421_p_dout0;
    output grp_sin_or_cos_double_s_fu_421_p_start;
    input grp_sin_or_cos_double_s_fu_421_p_ready;
    input grp_sin_or_cos_double_s_fu_421_p_done;
    input grp_sin_or_cos_double_s_fu_421_p_idle;
    output [63:0] grp_sin_or_cos_double_s_fu_432_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_432_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_432_p_dout0;
    output grp_sin_or_cos_double_s_fu_432_p_start;
    input grp_sin_or_cos_double_s_fu_432_p_ready;
    input grp_sin_or_cos_double_s_fu_432_p_done;
    input grp_sin_or_cos_double_s_fu_432_p_idle;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[16:0] pf_address0;
    reg pf_ce0;
    reg[31:0] pf_we0;
    reg[255:0] pf_d0;

    (* fsm_encoding = "none" *) reg   [242:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    reg   [30:0] seed;
    wire   [31:0] grp_fu_266_p2;
    reg   [31:0] reg_406;
    wire    ap_CS_fsm_state5;
    wire    ap_CS_fsm_state12;
    reg   [63:0] reg_411;
    wire    ap_CS_fsm_state7;
    wire    ap_CS_fsm_state79;
    wire    grp_atan2_cordic_double_s_fu_188_ap_done;
    wire    grp_sin_or_cos_double_s_fu_196_ap_done;
    wire    grp_sin_or_cos_double_s_fu_234_ap_done;
    reg    ap_block_state79_on_subcall_done;
    wire    ap_CS_fsm_state175;
    wire    ap_CS_fsm_state182;
    wire    ap_CS_fsm_state193;
    wire    ap_CS_fsm_state200;
    wire   [63:0] grp_fu_313_p1;
    reg   [63:0] reg_419;
    reg   [63:0] reg_427;
    wire    ap_CS_fsm_state14;
    wire    ap_CS_fsm_state21;
    wire    ap_CS_fsm_state36;
    wire    ap_CS_fsm_state93;
    reg   [63:0] reg_439;
    wire    ap_CS_fsm_state29;
    wire    ap_CS_fsm_state77;
    wire    ap_CS_fsm_state99;
    wire    ap_CS_fsm_state163;
    wire    ap_CS_fsm_state189;
    wire    ap_CS_fsm_state225;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_done;
    reg    ap_block_state225_on_subcall_done;
    wire    ap_CS_fsm_state232;
    reg   [63:0] reg_448;
    wire    ap_CS_fsm_state100;
    wire    ap_CS_fsm_state107;
    wire   [30:0] grp_fu_381_p2;
    reg   [30:0] reg_457;
    wire    ap_CS_fsm_state38;
    wire    ap_CS_fsm_state41;
    wire    ap_CS_fsm_state44;
    wire    ap_CS_fsm_state47;
    wire    ap_CS_fsm_state50;
    wire    ap_CS_fsm_state57;
    wire   [31:0] grp_fu_295_p1;
    reg   [31:0] reg_461;
    wire    ap_CS_fsm_state45;
    wire    ap_CS_fsm_state51;
    wire    ap_CS_fsm_state64;
    wire   [31:0] grp_fu_280_p2;
    reg   [31:0] reg_466;
    wire    ap_CS_fsm_state49;
    wire    ap_CS_fsm_state55;
    wire    ap_CS_fsm_state61;
    wire    ap_CS_fsm_state68;
    wire   [63:0] grp_fu_343_p2;
    reg   [63:0] reg_471;
    reg   [63:0] reg_478;
    wire    ap_CS_fsm_state218;
    reg   [63:0] reg_483;
    wire    ap_CS_fsm_state86;
    wire    ap_CS_fsm_state207;
    wire   [63:0] grp_fu_376_p2;
    reg   [63:0] reg_492;
    wire    ap_CS_fsm_state92;
    wire    ap_CS_fsm_state104;
    reg   [63:0] reg_497;
    wire    ap_CS_fsm_state235;
    reg   [63:0] reg_501;
    wire    ap_CS_fsm_state209;
    reg   [63:0] reg_505;
    wire    ap_CS_fsm_state114;
    wire    ap_CS_fsm_state169;
    wire   [63:0] grp_fu_349_p2;
    reg   [63:0] reg_512;
    wire   [63:0] grp_fu_353_p2;
    reg   [63:0] reg_518;
    reg   [63:0] reg_524;
    wire    ap_CS_fsm_state105;
    reg   [63:0] reg_530;
    wire    ap_CS_fsm_state196;
    wire    ap_CS_fsm_state216;
    wire    ap_CS_fsm_state242;
    reg   [63:0] reg_538;
    reg   [63:0] reg_545;
    wire    ap_CS_fsm_state121;
    wire    ap_CS_fsm_state223;
    reg   [63:0] reg_551;
    wire    ap_CS_fsm_state156;
    wire    ap_CS_fsm_state168;
    wire    ap_CS_fsm_state178;
    reg   [63:0] reg_557;
    wire    ap_CS_fsm_state162;
    wire    ap_CS_fsm_state171;
    wire   [31:0] grp_fu_304_p1;
    reg   [31:0] reg_563;
    wire    ap_CS_fsm_state173;
    wire    ap_CS_fsm_state180;
    wire    ap_CS_fsm_state191;
    wire    ap_CS_fsm_state198;
    wire   [31:0] grp_fu_307_p1;
    reg   [31:0] reg_568;
    wire  signed [30:0] grp_fu_573_p2;
    reg  signed [30:0] reg_579;
    wire    ap_CS_fsm_state39;
    wire    ap_CS_fsm_state42;
    reg  signed [30:0] reg_584;
    wire    ap_CS_fsm_state48;
    reg  signed [30:0] reg_589;
    wire    ap_CS_fsm_state58;
    wire   [31:0] grp_fu_272_p2;
    reg   [31:0] sub5_reg_889;
    wire    ap_CS_fsm_state8;
    wire   [63:0] bitcast_ln497_fu_610_p1;
    wire   [63:0] bitcast_ln497_1_fu_631_p1;
    reg   [63:0] thetaDiff_reg_915;
    wire   [63:0] bitcast_ln497_2_fu_651_p1;
    wire    ap_CS_fsm_state15;
    wire   [0:0] icmp_ln107_fu_674_p2;
    reg   [0:0] icmp_ln107_reg_926;
    wire    ap_CS_fsm_state22;
    wire   [0:0] icmp_ln107_1_fu_680_p2;
    reg   [0:0] icmp_ln107_1_reg_931;
    wire   [0:0] and_ln107_fu_690_p2;
    reg   [0:0] and_ln107_reg_936;
    wire    ap_CS_fsm_state23;
    wire   [31:0] zext_ln57_fu_706_p1;
    wire    ap_CS_fsm_state40;
    wire   [31:0] zext_ln57_2_fu_711_p1;
    wire    ap_CS_fsm_state46;
    reg   [63:0] conv2_i_reg_960;
    wire   [31:0] zext_ln57_4_fu_716_p1;
    wire    ap_CS_fsm_state52;
    reg   [63:0] conv2_i1_reg_970;
    wire   [31:0] zext_ln57_1_fu_727_p1;
    wire    ap_CS_fsm_state59;
    reg   [63:0] conv2_i2_reg_990;
    wire    ap_CS_fsm_state63;
    wire   [31:0] grp_fu_298_p1;
    reg   [31:0] conv1_i4_i1_reg_995;
    wire   [31:0] grp_fu_301_p1;
    reg   [31:0] conv1_i4_i2_reg_1000;
    wire   [31:0] grp_fu_285_p2;
    reg   [31:0] u2_1_reg_1005;
    wire   [31:0] grp_fu_290_p2;
    reg   [31:0] u2_2_reg_1010;
    reg   [63:0] conv3_i_reg_1015;
    wire    ap_CS_fsm_state70;
    reg   [63:0] conv3_i1_reg_1020;
    wire   [63:0] grp_fu_316_p1;
    reg   [63:0] conv3_i2_reg_1025;
    wire   [63:0] grp_atan2_cordic_double_s_fu_188_ap_return;
    reg   [63:0] tmp_s_reg_1030;
    reg   [63:0] tmp_18_reg_1035;
    wire   [63:0] grp_sin_or_cos_double_s_fu_234_ap_return;
    reg   [63:0] tmp_21_reg_1040;
    reg   [63:0] dTrans_reg_1050;
    wire   [63:0] trunc_ln116_fu_742_p1;
    reg   [63:0] trunc_ln116_reg_1057;
    reg   [63:0] trunc_ln117_1_reg_1062;
    wire   [63:0] bitcast_ln116_fu_756_p1;
    wire    ap_CS_fsm_state94;
    wire   [63:0] bitcast_ln116_1_fu_761_p1;
    wire   [63:0] bitcast_ln117_fu_766_p1;
    wire   [63:0] bitcast_ln117_1_fu_771_p1;
    reg   [63:0] bitcast_ln117_1_reg_1083;
    reg   [63:0] tmp_16_reg_1089;
    wire    ap_CS_fsm_state98;
    wire   [63:0] grp_fu_357_p2;
    reg   [63:0] mul13_reg_1094;
    reg   [63:0] mul_i2_reg_1099;
    wire    ap_CS_fsm_state111;
    wire   [63:0] grp_fu_327_p2;
    reg   [63:0] add6_reg_1104;
    wire   [63:0] grp_fu_371_p2;
    reg   [63:0] scaleH2_reg_1109;
    reg   [16:0] pf_addr_4_reg_1117;
    wire    ap_CS_fsm_state208;
    wire   [63:0] trunc_ln137_fu_800_p1;
    reg   [63:0] trunc_ln137_reg_1122;
    wire   [63:0] bitcast_ln135_fu_804_p1;
    wire    ap_CS_fsm_state210;
    wire   [63:0] bitcast_ln137_fu_809_p1;
    wire    ap_CS_fsm_state226;
    wire   [63:0] bitcast_ln138_fu_826_p1;
    wire    ap_CS_fsm_state236;
    wire    grp_atan2_cordic_double_s_fu_188_ap_start;
    wire    grp_atan2_cordic_double_s_fu_188_ap_idle;
    wire    grp_atan2_cordic_double_s_fu_188_ap_ready;
    wire   [63:0] grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din0;
    wire   [63:0] grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din1;
    wire   [0:0] grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_opcode;
    wire    grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_ce;
    wire   [63:0] grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din0;
    wire   [63:0] grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din1;
    wire   [4:0] grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_opcode;
    wire    grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_ce;
    wire    grp_sin_or_cos_double_s_fu_196_ap_ready;
    reg   [63:0] grp_sin_or_cos_double_s_fu_196_t_in;
    reg   [0:0] grp_sin_or_cos_double_s_fu_196_do_cos;
    wire    grp_sin_or_cos_double_s_fu_215_ap_ready;
    wire    grp_sin_or_cos_double_s_fu_234_ap_start;
    wire    grp_sin_or_cos_double_s_fu_234_ap_idle;
    wire    grp_sin_or_cos_double_s_fu_234_ap_ready;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_idle;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_ready;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_angle_assign_1_out;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_angle_assign_1_out_ap_vld;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din0;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din1;
    wire   [0:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_opcode;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_ce;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din0;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din1;
    wire   [4:0] grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_opcode;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_ce;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_idle;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_ready;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_angle_assign_3_out;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_angle_assign_3_out_ap_vld;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din0;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din1;
    wire   [0:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_opcode;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_ce;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din0;
    wire   [63:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din1;
    wire   [4:0] grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_opcode;
    wire    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_ce;
    reg    grp_atan2_cordic_double_s_fu_188_ap_start_reg;
    wire    ap_CS_fsm_state78;
    reg    grp_sin_or_cos_double_s_fu_196_ap_start_reg;
    wire    ap_CS_fsm_state217;
    wire    ap_CS_fsm_state224;
    reg    grp_sin_or_cos_double_s_fu_215_ap_start_reg;
    reg    grp_sin_or_cos_double_s_fu_234_ap_start_reg;
    reg    grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg;
    reg   [242:0] ap_NS_fsm;
    wire    ap_NS_fsm_state224;
    reg    grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg;
    wire    ap_CS_fsm_state227;
    wire   [63:0] zext_ln134_fu_790_p1;
    wire   [0:0] icmp_ln134_fu_778_p2;
    wire    ap_CS_fsm_state37;
    wire    ap_CS_fsm_state243;
    reg   [8:0] i_fu_126;
    wire   [8:0] add_ln134_fu_784_p2;
    wire    ap_CS_fsm_state24;
    wire    ap_CS_fsm_state233;
    wire   [255:0] zext_ln137_fu_821_p1;
    wire    ap_CS_fsm_state234;
    wire   [255:0] zext_ln139_fu_852_p1;
    reg   [31:0] grp_fu_266_p0;
    reg   [31:0] grp_fu_266_p1;
    wire    ap_CS_fsm_state65;
    reg   [31:0] grp_fu_295_p0;
    wire   [31:0] grp_fu_298_p0;
    wire   [31:0] grp_fu_301_p0;
    reg   [63:0] grp_fu_304_p0;
    wire    ap_CS_fsm_state172;
    wire    ap_CS_fsm_state179;
    wire    ap_CS_fsm_state190;
    wire    ap_CS_fsm_state197;
    reg   [63:0] grp_fu_307_p0;
    reg   [31:0] grp_fu_310_p0;
    wire    ap_CS_fsm_state6;
    wire    ap_CS_fsm_state13;
    wire    ap_CS_fsm_state56;
    wire    ap_CS_fsm_state62;
    wire    ap_CS_fsm_state69;
    wire    ap_CS_fsm_state174;
    wire    ap_CS_fsm_state181;
    wire    ap_CS_fsm_state192;
    wire    ap_CS_fsm_state199;
    reg   [31:0] grp_fu_313_p0;
    reg   [63:0] grp_fu_319_p0;
    reg   [63:0] grp_fu_319_p1;
    wire    ap_CS_fsm_state30;
    wire    ap_CS_fsm_state80;
    wire    ap_CS_fsm_state87;
    wire    ap_CS_fsm_state108;
    wire    ap_CS_fsm_state115;
    wire    ap_CS_fsm_state183;
    wire    ap_CS_fsm_state194;
    wire    ap_CS_fsm_state201;
    reg   [63:0] grp_fu_323_p0;
    reg   [63:0] grp_fu_323_p1;
    reg   [63:0] grp_fu_333_p0;
    reg   [63:0] grp_fu_333_p1;
    wire    ap_CS_fsm_state71;
    wire    ap_CS_fsm_state101;
    wire    ap_CS_fsm_state157;
    wire    ap_CS_fsm_state176;
    wire    ap_CS_fsm_state219;
    reg   [63:0] grp_fu_337_p0;
    reg   [63:0] grp_fu_337_p1;
    reg   [63:0] grp_fu_343_p0;
    reg   [63:0] grp_fu_343_p1;
    reg   [63:0] grp_fu_349_p0;
    reg   [63:0] grp_fu_353_p0;
    reg   [63:0] grp_fu_361_p0;
    reg   [63:0] grp_fu_361_p1;
    reg   [63:0] grp_fu_366_p1;
    wire    ap_CS_fsm_state106;
    wire    ap_CS_fsm_state112;
    wire    ap_CS_fsm_state122;
    reg   [63:0] grp_fu_376_p1;
    reg  signed [30:0] grp_fu_381_p0;
    wire    ap_CS_fsm_state43;
    wire   [63:0] data_fu_594_p1;
    wire   [62:0] trunc_ln479_fu_598_p1;
    wire   [63:0] t_fu_602_p3;
    wire   [63:0] data_1_fu_615_p1;
    wire   [62:0] trunc_ln479_1_fu_619_p1;
    wire   [63:0] t_1_fu_623_p3;
    wire   [63:0] data_2_fu_636_p1;
    wire   [62:0] trunc_ln479_2_fu_639_p1;
    wire   [63:0] t_2_fu_643_p3;
    wire   [63:0] bitcast_ln107_fu_656_p1;
    wire   [10:0] tmp_fu_660_p4;
    wire   [51:0] trunc_ln107_fu_670_p1;
    wire   [0:0] or_ln107_fu_686_p2;
    wire   [30:0] zext_ln57_5_fu_737_p0;
    wire   [63:0] bitcast_ln137_1_fu_817_p1;
    wire   [63:0] bitcast_ln46_fu_838_p1;
    wire   [63:0] bitcast_ln138_1_fu_831_p1;
    wire   [191:0] or_ln139_7_fu_842_p4;
    reg    grp_fu_310_ce;
    reg   [1:0] grp_fu_319_opcode;
    reg    grp_fu_319_ce;
    wire    ap_CS_fsm_state9;
    wire    ap_CS_fsm_state10;
    wire    ap_CS_fsm_state11;
    wire    ap_CS_fsm_state16;
    wire    ap_CS_fsm_state17;
    wire    ap_CS_fsm_state18;
    wire    ap_CS_fsm_state19;
    wire    ap_CS_fsm_state20;
    wire    ap_CS_fsm_state31;
    wire    ap_CS_fsm_state32;
    wire    ap_CS_fsm_state33;
    wire    ap_CS_fsm_state34;
    wire    ap_CS_fsm_state35;
    wire    ap_CS_fsm_state81;
    wire    ap_CS_fsm_state82;
    wire    ap_CS_fsm_state83;
    wire    ap_CS_fsm_state84;
    wire    ap_CS_fsm_state85;
    wire    ap_CS_fsm_state88;
    wire    ap_CS_fsm_state89;
    wire    ap_CS_fsm_state90;
    wire    ap_CS_fsm_state91;
    wire    ap_CS_fsm_state109;
    wire    ap_CS_fsm_state110;
    wire    ap_CS_fsm_state113;
    wire    ap_CS_fsm_state116;
    wire    ap_CS_fsm_state117;
    wire    ap_CS_fsm_state118;
    wire    ap_CS_fsm_state119;
    wire    ap_CS_fsm_state120;
    wire    ap_CS_fsm_state184;
    wire    ap_CS_fsm_state185;
    wire    ap_CS_fsm_state186;
    wire    ap_CS_fsm_state187;
    wire    ap_CS_fsm_state188;
    wire    ap_CS_fsm_state195;
    wire    ap_CS_fsm_state202;
    wire    ap_CS_fsm_state203;
    wire    ap_CS_fsm_state204;
    wire    ap_CS_fsm_state205;
    wire    ap_CS_fsm_state206;
    wire    ap_CS_fsm_state211;
    wire    ap_CS_fsm_state212;
    wire    ap_CS_fsm_state213;
    wire    ap_CS_fsm_state214;
    wire    ap_CS_fsm_state215;
    wire    ap_CS_fsm_state220;
    wire    ap_CS_fsm_state221;
    wire    ap_CS_fsm_state222;
    wire    ap_CS_fsm_state228;
    wire    ap_CS_fsm_state229;
    wire    ap_CS_fsm_state230;
    wire    ap_CS_fsm_state231;
    wire    ap_CS_fsm_state237;
    wire    ap_CS_fsm_state238;
    wire    ap_CS_fsm_state239;
    wire    ap_CS_fsm_state240;
    wire    ap_CS_fsm_state241;
    reg   [1:0] grp_fu_323_opcode;
    reg    grp_fu_323_ce;
    reg    grp_fu_333_ce;
    wire    ap_CS_fsm_state25;
    wire    ap_CS_fsm_state26;
    wire    ap_CS_fsm_state27;
    wire    ap_CS_fsm_state28;
    wire    ap_CS_fsm_state72;
    wire    ap_CS_fsm_state73;
    wire    ap_CS_fsm_state74;
    wire    ap_CS_fsm_state75;
    wire    ap_CS_fsm_state76;
    wire    ap_CS_fsm_state95;
    wire    ap_CS_fsm_state96;
    wire    ap_CS_fsm_state97;
    wire    ap_CS_fsm_state102;
    wire    ap_CS_fsm_state103;
    wire    ap_CS_fsm_state158;
    wire    ap_CS_fsm_state159;
    wire    ap_CS_fsm_state160;
    wire    ap_CS_fsm_state161;
    wire    ap_CS_fsm_state164;
    wire    ap_CS_fsm_state165;
    wire    ap_CS_fsm_state166;
    wire    ap_CS_fsm_state167;
    wire    ap_CS_fsm_state170;
    wire    ap_CS_fsm_state177;
    reg    grp_fu_361_ce;
    reg   [4:0] grp_fu_361_opcode;
    reg    grp_fu_366_ce;
    wire    ap_CS_fsm_state53;
    wire    ap_CS_fsm_state54;
    wire    ap_CS_fsm_state60;
    wire    ap_CS_fsm_state66;
    wire    ap_CS_fsm_state67;
    wire    ap_CS_fsm_state2;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    reg    grp_fu_376_ce;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_ST_fsm_state62_blk;
    wire    ap_ST_fsm_state63_blk;
    wire    ap_ST_fsm_state64_blk;
    wire    ap_ST_fsm_state65_blk;
    wire    ap_ST_fsm_state66_blk;
    wire    ap_ST_fsm_state67_blk;
    wire    ap_ST_fsm_state68_blk;
    wire    ap_ST_fsm_state69_blk;
    wire    ap_ST_fsm_state70_blk;
    wire    ap_ST_fsm_state71_blk;
    wire    ap_ST_fsm_state72_blk;
    wire    ap_ST_fsm_state73_blk;
    wire    ap_ST_fsm_state74_blk;
    wire    ap_ST_fsm_state75_blk;
    wire    ap_ST_fsm_state76_blk;
    wire    ap_ST_fsm_state77_blk;
    wire    ap_ST_fsm_state78_blk;
    reg    ap_ST_fsm_state79_blk;
    wire    ap_ST_fsm_state80_blk;
    wire    ap_ST_fsm_state81_blk;
    wire    ap_ST_fsm_state82_blk;
    wire    ap_ST_fsm_state83_blk;
    wire    ap_ST_fsm_state84_blk;
    wire    ap_ST_fsm_state85_blk;
    wire    ap_ST_fsm_state86_blk;
    wire    ap_ST_fsm_state87_blk;
    wire    ap_ST_fsm_state88_blk;
    wire    ap_ST_fsm_state89_blk;
    wire    ap_ST_fsm_state90_blk;
    wire    ap_ST_fsm_state91_blk;
    wire    ap_ST_fsm_state92_blk;
    wire    ap_ST_fsm_state93_blk;
    wire    ap_ST_fsm_state94_blk;
    wire    ap_ST_fsm_state95_blk;
    wire    ap_ST_fsm_state96_blk;
    wire    ap_ST_fsm_state97_blk;
    wire    ap_ST_fsm_state98_blk;
    wire    ap_ST_fsm_state99_blk;
    wire    ap_ST_fsm_state100_blk;
    wire    ap_ST_fsm_state101_blk;
    wire    ap_ST_fsm_state102_blk;
    wire    ap_ST_fsm_state103_blk;
    wire    ap_ST_fsm_state104_blk;
    wire    ap_ST_fsm_state105_blk;
    wire    ap_ST_fsm_state106_blk;
    wire    ap_ST_fsm_state107_blk;
    wire    ap_ST_fsm_state108_blk;
    wire    ap_ST_fsm_state109_blk;
    wire    ap_ST_fsm_state110_blk;
    wire    ap_ST_fsm_state111_blk;
    wire    ap_ST_fsm_state112_blk;
    wire    ap_ST_fsm_state113_blk;
    wire    ap_ST_fsm_state114_blk;
    wire    ap_ST_fsm_state115_blk;
    wire    ap_ST_fsm_state116_blk;
    wire    ap_ST_fsm_state117_blk;
    wire    ap_ST_fsm_state118_blk;
    wire    ap_ST_fsm_state119_blk;
    wire    ap_ST_fsm_state120_blk;
    wire    ap_ST_fsm_state121_blk;
    wire    ap_ST_fsm_state122_blk;
    wire    ap_ST_fsm_state123_blk;
    wire    ap_ST_fsm_state124_blk;
    wire    ap_ST_fsm_state125_blk;
    wire    ap_ST_fsm_state126_blk;
    wire    ap_ST_fsm_state127_blk;
    wire    ap_ST_fsm_state128_blk;
    wire    ap_ST_fsm_state129_blk;
    wire    ap_ST_fsm_state130_blk;
    wire    ap_ST_fsm_state131_blk;
    wire    ap_ST_fsm_state132_blk;
    wire    ap_ST_fsm_state133_blk;
    wire    ap_ST_fsm_state134_blk;
    wire    ap_ST_fsm_state135_blk;
    wire    ap_ST_fsm_state136_blk;
    wire    ap_ST_fsm_state137_blk;
    wire    ap_ST_fsm_state138_blk;
    wire    ap_ST_fsm_state139_blk;
    wire    ap_ST_fsm_state140_blk;
    wire    ap_ST_fsm_state141_blk;
    wire    ap_ST_fsm_state142_blk;
    wire    ap_ST_fsm_state143_blk;
    wire    ap_ST_fsm_state144_blk;
    wire    ap_ST_fsm_state145_blk;
    wire    ap_ST_fsm_state146_blk;
    wire    ap_ST_fsm_state147_blk;
    wire    ap_ST_fsm_state148_blk;
    wire    ap_ST_fsm_state149_blk;
    wire    ap_ST_fsm_state150_blk;
    wire    ap_ST_fsm_state151_blk;
    wire    ap_ST_fsm_state152_blk;
    wire    ap_ST_fsm_state153_blk;
    wire    ap_ST_fsm_state154_blk;
    wire    ap_ST_fsm_state155_blk;
    wire    ap_ST_fsm_state156_blk;
    wire    ap_ST_fsm_state157_blk;
    wire    ap_ST_fsm_state158_blk;
    wire    ap_ST_fsm_state159_blk;
    wire    ap_ST_fsm_state160_blk;
    wire    ap_ST_fsm_state161_blk;
    wire    ap_ST_fsm_state162_blk;
    wire    ap_ST_fsm_state163_blk;
    wire    ap_ST_fsm_state164_blk;
    wire    ap_ST_fsm_state165_blk;
    wire    ap_ST_fsm_state166_blk;
    wire    ap_ST_fsm_state167_blk;
    wire    ap_ST_fsm_state168_blk;
    wire    ap_ST_fsm_state169_blk;
    wire    ap_ST_fsm_state170_blk;
    wire    ap_ST_fsm_state171_blk;
    wire    ap_ST_fsm_state172_blk;
    wire    ap_ST_fsm_state173_blk;
    wire    ap_ST_fsm_state174_blk;
    wire    ap_ST_fsm_state175_blk;
    wire    ap_ST_fsm_state176_blk;
    wire    ap_ST_fsm_state177_blk;
    wire    ap_ST_fsm_state178_blk;
    wire    ap_ST_fsm_state179_blk;
    wire    ap_ST_fsm_state180_blk;
    wire    ap_ST_fsm_state181_blk;
    wire    ap_ST_fsm_state182_blk;
    wire    ap_ST_fsm_state183_blk;
    wire    ap_ST_fsm_state184_blk;
    wire    ap_ST_fsm_state185_blk;
    wire    ap_ST_fsm_state186_blk;
    wire    ap_ST_fsm_state187_blk;
    wire    ap_ST_fsm_state188_blk;
    wire    ap_ST_fsm_state189_blk;
    wire    ap_ST_fsm_state190_blk;
    wire    ap_ST_fsm_state191_blk;
    wire    ap_ST_fsm_state192_blk;
    wire    ap_ST_fsm_state193_blk;
    wire    ap_ST_fsm_state194_blk;
    wire    ap_ST_fsm_state195_blk;
    wire    ap_ST_fsm_state196_blk;
    wire    ap_ST_fsm_state197_blk;
    wire    ap_ST_fsm_state198_blk;
    wire    ap_ST_fsm_state199_blk;
    wire    ap_ST_fsm_state200_blk;
    wire    ap_ST_fsm_state201_blk;
    wire    ap_ST_fsm_state202_blk;
    wire    ap_ST_fsm_state203_blk;
    wire    ap_ST_fsm_state204_blk;
    wire    ap_ST_fsm_state205_blk;
    wire    ap_ST_fsm_state206_blk;
    wire    ap_ST_fsm_state207_blk;
    wire    ap_ST_fsm_state208_blk;
    wire    ap_ST_fsm_state209_blk;
    wire    ap_ST_fsm_state210_blk;
    wire    ap_ST_fsm_state211_blk;
    wire    ap_ST_fsm_state212_blk;
    wire    ap_ST_fsm_state213_blk;
    wire    ap_ST_fsm_state214_blk;
    wire    ap_ST_fsm_state215_blk;
    wire    ap_ST_fsm_state216_blk;
    wire    ap_ST_fsm_state217_blk;
    reg    ap_ST_fsm_state218_blk;
    wire    ap_ST_fsm_state219_blk;
    wire    ap_ST_fsm_state220_blk;
    wire    ap_ST_fsm_state221_blk;
    wire    ap_ST_fsm_state222_blk;
    wire    ap_ST_fsm_state223_blk;
    wire    ap_ST_fsm_state224_blk;
    reg    ap_ST_fsm_state225_blk;
    wire    ap_ST_fsm_state226_blk;
    reg    ap_ST_fsm_state227_blk;
    wire    ap_ST_fsm_state228_blk;
    wire    ap_ST_fsm_state229_blk;
    wire    ap_ST_fsm_state230_blk;
    wire    ap_ST_fsm_state231_blk;
    wire    ap_ST_fsm_state232_blk;
    wire    ap_ST_fsm_state233_blk;
    wire    ap_ST_fsm_state234_blk;
    wire    ap_ST_fsm_state235_blk;
    wire    ap_ST_fsm_state236_blk;
    wire    ap_ST_fsm_state237_blk;
    wire    ap_ST_fsm_state238_blk;
    wire    ap_ST_fsm_state239_blk;
    wire    ap_ST_fsm_state240_blk;
    wire    ap_ST_fsm_state241_blk;
    wire    ap_ST_fsm_state242_blk;
    wire    ap_ST_fsm_state243_blk;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 243'd1;
        #0 seed = 31'd123456789;
        #0 grp_atan2_cordic_double_s_fu_188_ap_start_reg = 1'b0;
        #0 grp_sin_or_cos_double_s_fu_196_ap_start_reg = 1'b0;
        #0 grp_sin_or_cos_double_s_fu_215_ap_start_reg = 1'b0;
        #0 grp_sin_or_cos_double_s_fu_234_ap_start_reg = 1'b0;
        #0 grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg = 1'b0;
        #0 grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg = 1'b0;
        #0 i_fu_126 = 9'd0;
    end

    main_atan2_cordic_double_s grp_atan2_cordic_double_s_fu_188 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_atan2_cordic_double_s_fu_188_ap_start),
        .ap_done(grp_atan2_cordic_double_s_fu_188_ap_done),
        .ap_idle(grp_atan2_cordic_double_s_fu_188_ap_idle),
        .ap_ready(grp_atan2_cordic_double_s_fu_188_ap_ready),
        .y_in(reg_419),
        .x_in(reg_411),
        .ap_return(grp_atan2_cordic_double_s_fu_188_ap_return),
        .grp_fu_323_p_din0(grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din0),
        .grp_fu_323_p_din1(grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din1),
        .grp_fu_323_p_opcode(grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_opcode),
        .grp_fu_323_p_dout0(grp_fu_401_p_dout0),
        .grp_fu_323_p_ce(grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_ce),
        .grp_fu_361_p_din0(grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din0),
        .grp_fu_361_p_din1(grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din1),
        .grp_fu_361_p_opcode(grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_opcode),
        .grp_fu_361_p_dout0(grp_fu_413_p_dout0),
        .grp_fu_361_p_ce(grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_ce)
    );

    main_sin_or_cos_double_s grp_sin_or_cos_double_s_fu_234 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_sin_or_cos_double_s_fu_234_ap_start),
        .ap_done(grp_sin_or_cos_double_s_fu_234_ap_done),
        .ap_idle(grp_sin_or_cos_double_s_fu_234_ap_idle),
        .ap_ready(grp_sin_or_cos_double_s_fu_234_ap_ready),
        .t_in(reg_471),
        .do_cos(1'd1),
        .ap_return(grp_sin_or_cos_double_s_fu_234_ap_return)
    );

    main_updateMotion_Pipeline_VITIS_LOOP_45_1 grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start),
        .ap_done(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_done),
        .ap_idle(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_idle),
        .ap_ready(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_ready),
        .angle_assign(reg_545),
        .angle_assign_1_out(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_angle_assign_1_out),
        .angle_assign_1_out_ap_vld(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_angle_assign_1_out_ap_vld),
        .grp_fu_323_p_din0(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din0),
        .grp_fu_323_p_din1(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din1),
        .grp_fu_323_p_opcode(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_opcode),
        .grp_fu_323_p_dout0(grp_fu_401_p_dout0),
        .grp_fu_323_p_ce(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_ce),
        .grp_fu_361_p_din0(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din0),
        .grp_fu_361_p_din1(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din1),
        .grp_fu_361_p_opcode(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_opcode),
        .grp_fu_361_p_dout0(grp_fu_413_p_dout0),
        .grp_fu_361_p_ce(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_ce)
    );

    main_updateMotion_Pipeline_VITIS_LOOP_46_2 grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start),
        .ap_done(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done),
        .ap_idle(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_idle),
        .ap_ready(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_ready),
        .angle_assign_1_reload(grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_angle_assign_1_out),
        .angle_assign_3_out(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_angle_assign_3_out),
        .angle_assign_3_out_ap_vld(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_angle_assign_3_out_ap_vld),
        .grp_fu_323_p_din0(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din0),
        .grp_fu_323_p_din1(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din1),
        .grp_fu_323_p_opcode(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_opcode),
        .grp_fu_323_p_dout0(grp_fu_401_p_dout0),
        .grp_fu_323_p_ce(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_ce),
        .grp_fu_361_p_din0(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din0),
        .grp_fu_361_p_din1(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din1),
        .grp_fu_361_p_opcode(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_opcode),
        .grp_fu_361_p_dout0(grp_fu_413_p_dout0),
        .grp_fu_361_p_ce(grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_ce)
    );

    main_fsub_32ns_32ns_32_5_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fsub_32ns_32ns_32_5_full_dsp_1_U92 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_266_p0),
        .din1(grp_fu_266_p1),
        .ce(1'b1),
        .dout(grp_fu_266_p2)
    );

    main_fsub_32ns_32ns_32_5_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fsub_32ns_32ns_32_5_full_dsp_1_U93 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(currOdometry_0_1_val),
        .din1(prevOdometry_0_1_val),
        .ce(1'b1),
        .dout(grp_fu_272_p2)
    );

    main_fmul_32ns_32ns_32_4_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fmul_32ns_32ns_32_4_max_dsp_1_U94 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(reg_461),
        .din1(32'd805306368),
        .ce(1'b1),
        .dout(grp_fu_280_p2)
    );

    main_fmul_32ns_32ns_32_4_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fmul_32ns_32ns_32_4_max_dsp_1_U95 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(conv1_i4_i1_reg_995),
        .din1(32'd805306368),
        .ce(1'b1),
        .dout(grp_fu_285_p2)
    );

    main_fmul_32ns_32ns_32_4_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fmul_32ns_32ns_32_4_max_dsp_1_U96 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(conv1_i4_i2_reg_1000),
        .din1(32'd805306368),
        .ce(1'b1),
        .dout(grp_fu_290_p2)
    );

    main_uitofp_32ns_32_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(32)
    ) uitofp_32ns_32_6_no_dsp_1_U97 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_295_p0),
        .ce(1'b1),
        .dout(grp_fu_295_p1)
    );

    main_uitofp_32ns_32_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(32)
    ) uitofp_32ns_32_6_no_dsp_1_U98 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_298_p0),
        .ce(1'b1),
        .dout(grp_fu_298_p1)
    );

    main_uitofp_32ns_32_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(32)
    ) uitofp_32ns_32_6_no_dsp_1_U99 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_301_p0),
        .ce(1'b1),
        .dout(grp_fu_301_p1)
    );

    main_fptrunc_64ns_32_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .dout_WIDTH(32)
    ) fptrunc_64ns_32_2_no_dsp_1_U100 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_304_p0),
        .ce(1'b1),
        .dout(grp_fu_304_p1)
    );

    main_fptrunc_64ns_32_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .dout_WIDTH(32)
    ) fptrunc_64ns_32_2_no_dsp_1_U101 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_307_p0),
        .ce(1'b1),
        .dout(grp_fu_307_p1)
    );

    main_fpext_32ns_64_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) fpext_32ns_64_2_no_dsp_1_U103 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_313_p0),
        .ce(1'b1),
        .dout(grp_fu_313_p1)
    );

    main_fpext_32ns_64_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) fpext_32ns_64_2_no_dsp_1_U104 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(u2_2_reg_1010),
        .ce(1'b1),
        .dout(grp_fu_316_p1)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U107 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul13_reg_1094),
        .din1(reg_448),
        .ce(1'b1),
        .dout(grp_fu_327_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U110 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_343_p0),
        .din1(grp_fu_343_p1),
        .ce(1'b1),
        .dout(grp_fu_343_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U111 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_349_p0),
        .din1(reg_483),
        .ce(1'b1),
        .dout(grp_fu_349_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U112 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_353_p0),
        .din1(reg_427),
        .ce(1'b1),
        .dout(grp_fu_353_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U113 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(reg_518),
        .din1(reg_427),
        .ce(1'b1),
        .dout(grp_fu_357_p2)
    );

    main_dsqrt_64ns_64ns_64_57_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(57),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsqrt_64ns_64ns_64_57_no_dsp_1_U116 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd0),
        .din1(add6_reg_1104),
        .ce(1'b1),
        .dout(grp_fu_371_p2)
    );

    main_dlog_64ns_64ns_64_41_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(41),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dlog_64ns_64ns_64_41_full_dsp_1_U117 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd0),
        .din1(grp_fu_376_p1),
        .ce(grp_fu_376_ce),
        .dout(grp_fu_376_p2)
    );

    main_mul_31s_31s_31_2_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(31),
        .din1_WIDTH(31),
        .dout_WIDTH(31)
    ) mul_31s_31s_31_2_1_U118 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_381_p0),
        .din1(31'd1103515245),
        .ce(1'b1),
        .dout(grp_fu_381_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_atan2_cordic_double_s_fu_188_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state78)) begin
                grp_atan2_cordic_double_s_fu_188_ap_start_reg <= 1'b1;
            end else if ((grp_atan2_cordic_double_s_fu_188_ap_ready == 1'b1)) begin
                grp_atan2_cordic_double_s_fu_188_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_196_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state217) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state224))) begin
                grp_sin_or_cos_double_s_fu_196_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_196_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_196_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_215_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state78)) begin
                grp_sin_or_cos_double_s_fu_215_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_215_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_215_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_sin_or_cos_double_s_fu_234_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state78)) begin
                grp_sin_or_cos_double_s_fu_234_ap_start_reg <= 1'b1;
            end else if ((grp_sin_or_cos_double_s_fu_234_ap_ready == 1'b1)) begin
                grp_sin_or_cos_double_s_fu_234_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state223) & (1'b1 == ap_NS_fsm_state224))) begin
                grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg <= 1'b1;
            end else if ((grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_ready == 1'b1)) begin
                grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state226)) begin
                grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg <= 1'b1;
            end else if ((grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_ready == 1'b1)) begin
                grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state24)) begin
            i_fu_126 <= 9'd0;
        end else if (((1'b1 == ap_CS_fsm_state208) & (icmp_ln134_fu_778_p2 == 1'd0) & (1'd0 == and_ln107_reg_936))) begin
            i_fu_126 <= add_ln134_fu_784_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state114)) begin
            add6_reg_1104 <= grp_fu_327_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state23)) begin
            and_ln107_reg_936 <= and_ln107_fu_690_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state94)) begin
            bitcast_ln117_1_reg_1083 <= bitcast_ln117_1_fu_771_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state64)) begin
            conv1_i4_i1_reg_995  <= grp_fu_298_p1;
            conv1_i4_i2_reg_1000 <= grp_fu_301_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state57)) begin
            conv2_i1_reg_970 <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state63)) begin
            conv2_i2_reg_990 <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state51)) begin
            conv2_i_reg_960 <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state70)) begin
            conv3_i1_reg_1020 <= grp_fu_313_p1;
            conv3_i2_reg_1025 <= grp_fu_316_p1;
            conv3_i_reg_1015  <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state93)) begin
            dTrans_reg_1050 <= grp_fu_417_p_dout0;
            trunc_ln116_reg_1057 <= trunc_ln116_fu_742_p1;
            trunc_ln117_1_reg_1062 <= {{pf_q0[255:192]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state22)) begin
            icmp_ln107_1_reg_931 <= icmp_ln107_1_fu_680_p2;
            icmp_ln107_reg_926   <= icmp_ln107_fu_674_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state107)) begin
            mul13_reg_1094 <= grp_fu_357_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state111)) begin
            mul_i2_reg_1099 <= grp_fu_405_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state208)) begin
            pf_addr_4_reg_1117[8 : 0] <= zext_ln134_fu_790_p1[8 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5))) begin
            reg_406 <= grp_fu_266_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state200) | (1'b1 == ap_CS_fsm_state193) | (1'b1 == ap_CS_fsm_state182) | (1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state7) | ((1'b0 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79)))) begin
            reg_411 <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state193) | (1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state7))) begin
            reg_419 <= grp_fu_313_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state93) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state200))) begin
            reg_427 <= grp_fu_397_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state232) | (1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state163) | (1'b1 == ap_CS_fsm_state99) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state182) | ((1'b0 == ap_block_state225_on_subcall_done) & (1'b1 == ap_CS_fsm_state225)))) begin
            reg_439 <= grp_fu_405_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state107) | (1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state182))) begin
            reg_448 <= grp_fu_409_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state41) | (1'b1 == ap_CS_fsm_state38))) begin
            reg_457 <= grp_fu_381_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state45) | (1'b1 == ap_CS_fsm_state57))) begin
            reg_461 <= grp_fu_295_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state49))) begin
            reg_466 <= grp_fu_280_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state107) | (1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state77))) begin
            reg_471 <= grp_fu_343_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((grp_sin_or_cos_double_s_fu_196_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state218)) | ((1'b0 == ap_block_state225_on_subcall_done) & (1'b1 == ap_CS_fsm_state225)) | ((1'b0 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79)))) begin
            reg_478 <= grp_sin_or_cos_double_s_fu_421_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state207) | (1'b1 == ap_CS_fsm_state86))) begin
            reg_483 <= grp_fu_397_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state104) | (1'b1 == ap_CS_fsm_state92))) begin
            reg_492 <= grp_fu_376_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state235) | (1'b1 == ap_CS_fsm_state93))) begin
            reg_497 <= {{pf_q0[127:64]}};
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state209) | (1'b1 == ap_CS_fsm_state93))) begin
            reg_501 <= {{pf_q0[191:128]}};
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state169) | (1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state107) | (1'b1 == ap_CS_fsm_state100))) begin
            reg_505 <= grp_fu_405_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state107) | (1'b1 == ap_CS_fsm_state100))) begin
            reg_512 <= grp_fu_349_p2;
            reg_518 <= grp_fu_353_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state105) | (1'b1 == ap_CS_fsm_state175))) begin
            reg_524 <= grp_fu_405_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state242) | (1'b1 == ap_CS_fsm_state216) | (1'b1 == ap_CS_fsm_state196) | (1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state232) | (1'b1 == ap_CS_fsm_state189))) begin
            reg_530 <= grp_fu_397_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state200))) begin
            reg_538 <= grp_fu_401_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state223) | (1'b1 == ap_CS_fsm_state121))) begin
            reg_545 <= grp_fu_397_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state178) | (1'b1 == ap_CS_fsm_state168) | (1'b1 == ap_CS_fsm_state156))) begin
            reg_551 <= grp_fu_417_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state171) | (1'b1 == ap_CS_fsm_state162))) begin
            reg_557 <= grp_fu_417_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state198) | (1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state180) | (1'b1 == ap_CS_fsm_state173))) begin
            reg_563 <= grp_fu_304_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state173))) begin
            reg_568 <= grp_fu_307_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state42) | (1'b1 == ap_CS_fsm_state39))) begin
            reg_579 <= grp_fu_573_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state45))) begin
            reg_584 <= grp_fu_573_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state51))) begin
            reg_589 <= grp_fu_573_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state171)) begin
            scaleH2_reg_1109 <= grp_fu_371_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state58)) begin
            seed <= grp_fu_573_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            sub5_reg_889 <= grp_fu_272_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state14)) begin
            thetaDiff_reg_915 <= grp_fu_394_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state98)) begin
            tmp_16_reg_1089 <= grp_fu_376_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state79)) begin
            tmp_18_reg_1035 <= grp_sin_or_cos_double_s_fu_432_p_dout0;
            tmp_21_reg_1040 <= grp_sin_or_cos_double_s_fu_234_ap_return;
            tmp_s_reg_1030  <= grp_atan2_cordic_double_s_fu_188_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            trunc_ln137_reg_1122 <= trunc_ln137_fu_800_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state68)) begin
            u2_1_reg_1005 <= grp_fu_285_p2;
            u2_2_reg_1010 <= grp_fu_290_p2;
        end
    end

    assign ap_ST_fsm_state100_blk = 1'b0;

    assign ap_ST_fsm_state101_blk = 1'b0;

    assign ap_ST_fsm_state102_blk = 1'b0;

    assign ap_ST_fsm_state103_blk = 1'b0;

    assign ap_ST_fsm_state104_blk = 1'b0;

    assign ap_ST_fsm_state105_blk = 1'b0;

    assign ap_ST_fsm_state106_blk = 1'b0;

    assign ap_ST_fsm_state107_blk = 1'b0;

    assign ap_ST_fsm_state108_blk = 1'b0;

    assign ap_ST_fsm_state109_blk = 1'b0;

    assign ap_ST_fsm_state10_blk  = 1'b0;

    assign ap_ST_fsm_state110_blk = 1'b0;

    assign ap_ST_fsm_state111_blk = 1'b0;

    assign ap_ST_fsm_state112_blk = 1'b0;

    assign ap_ST_fsm_state113_blk = 1'b0;

    assign ap_ST_fsm_state114_blk = 1'b0;

    assign ap_ST_fsm_state115_blk = 1'b0;

    assign ap_ST_fsm_state116_blk = 1'b0;

    assign ap_ST_fsm_state117_blk = 1'b0;

    assign ap_ST_fsm_state118_blk = 1'b0;

    assign ap_ST_fsm_state119_blk = 1'b0;

    assign ap_ST_fsm_state11_blk  = 1'b0;

    assign ap_ST_fsm_state120_blk = 1'b0;

    assign ap_ST_fsm_state121_blk = 1'b0;

    assign ap_ST_fsm_state122_blk = 1'b0;

    assign ap_ST_fsm_state123_blk = 1'b0;

    assign ap_ST_fsm_state124_blk = 1'b0;

    assign ap_ST_fsm_state125_blk = 1'b0;

    assign ap_ST_fsm_state126_blk = 1'b0;

    assign ap_ST_fsm_state127_blk = 1'b0;

    assign ap_ST_fsm_state128_blk = 1'b0;

    assign ap_ST_fsm_state129_blk = 1'b0;

    assign ap_ST_fsm_state12_blk  = 1'b0;

    assign ap_ST_fsm_state130_blk = 1'b0;

    assign ap_ST_fsm_state131_blk = 1'b0;

    assign ap_ST_fsm_state132_blk = 1'b0;

    assign ap_ST_fsm_state133_blk = 1'b0;

    assign ap_ST_fsm_state134_blk = 1'b0;

    assign ap_ST_fsm_state135_blk = 1'b0;

    assign ap_ST_fsm_state136_blk = 1'b0;

    assign ap_ST_fsm_state137_blk = 1'b0;

    assign ap_ST_fsm_state138_blk = 1'b0;

    assign ap_ST_fsm_state139_blk = 1'b0;

    assign ap_ST_fsm_state13_blk  = 1'b0;

    assign ap_ST_fsm_state140_blk = 1'b0;

    assign ap_ST_fsm_state141_blk = 1'b0;

    assign ap_ST_fsm_state142_blk = 1'b0;

    assign ap_ST_fsm_state143_blk = 1'b0;

    assign ap_ST_fsm_state144_blk = 1'b0;

    assign ap_ST_fsm_state145_blk = 1'b0;

    assign ap_ST_fsm_state146_blk = 1'b0;

    assign ap_ST_fsm_state147_blk = 1'b0;

    assign ap_ST_fsm_state148_blk = 1'b0;

    assign ap_ST_fsm_state149_blk = 1'b0;

    assign ap_ST_fsm_state14_blk  = 1'b0;

    assign ap_ST_fsm_state150_blk = 1'b0;

    assign ap_ST_fsm_state151_blk = 1'b0;

    assign ap_ST_fsm_state152_blk = 1'b0;

    assign ap_ST_fsm_state153_blk = 1'b0;

    assign ap_ST_fsm_state154_blk = 1'b0;

    assign ap_ST_fsm_state155_blk = 1'b0;

    assign ap_ST_fsm_state156_blk = 1'b0;

    assign ap_ST_fsm_state157_blk = 1'b0;

    assign ap_ST_fsm_state158_blk = 1'b0;

    assign ap_ST_fsm_state159_blk = 1'b0;

    assign ap_ST_fsm_state15_blk  = 1'b0;

    assign ap_ST_fsm_state160_blk = 1'b0;

    assign ap_ST_fsm_state161_blk = 1'b0;

    assign ap_ST_fsm_state162_blk = 1'b0;

    assign ap_ST_fsm_state163_blk = 1'b0;

    assign ap_ST_fsm_state164_blk = 1'b0;

    assign ap_ST_fsm_state165_blk = 1'b0;

    assign ap_ST_fsm_state166_blk = 1'b0;

    assign ap_ST_fsm_state167_blk = 1'b0;

    assign ap_ST_fsm_state168_blk = 1'b0;

    assign ap_ST_fsm_state169_blk = 1'b0;

    assign ap_ST_fsm_state16_blk  = 1'b0;

    assign ap_ST_fsm_state170_blk = 1'b0;

    assign ap_ST_fsm_state171_blk = 1'b0;

    assign ap_ST_fsm_state172_blk = 1'b0;

    assign ap_ST_fsm_state173_blk = 1'b0;

    assign ap_ST_fsm_state174_blk = 1'b0;

    assign ap_ST_fsm_state175_blk = 1'b0;

    assign ap_ST_fsm_state176_blk = 1'b0;

    assign ap_ST_fsm_state177_blk = 1'b0;

    assign ap_ST_fsm_state178_blk = 1'b0;

    assign ap_ST_fsm_state179_blk = 1'b0;

    assign ap_ST_fsm_state17_blk  = 1'b0;

    assign ap_ST_fsm_state180_blk = 1'b0;

    assign ap_ST_fsm_state181_blk = 1'b0;

    assign ap_ST_fsm_state182_blk = 1'b0;

    assign ap_ST_fsm_state183_blk = 1'b0;

    assign ap_ST_fsm_state184_blk = 1'b0;

    assign ap_ST_fsm_state185_blk = 1'b0;

    assign ap_ST_fsm_state186_blk = 1'b0;

    assign ap_ST_fsm_state187_blk = 1'b0;

    assign ap_ST_fsm_state188_blk = 1'b0;

    assign ap_ST_fsm_state189_blk = 1'b0;

    assign ap_ST_fsm_state18_blk  = 1'b0;

    assign ap_ST_fsm_state190_blk = 1'b0;

    assign ap_ST_fsm_state191_blk = 1'b0;

    assign ap_ST_fsm_state192_blk = 1'b0;

    assign ap_ST_fsm_state193_blk = 1'b0;

    assign ap_ST_fsm_state194_blk = 1'b0;

    assign ap_ST_fsm_state195_blk = 1'b0;

    assign ap_ST_fsm_state196_blk = 1'b0;

    assign ap_ST_fsm_state197_blk = 1'b0;

    assign ap_ST_fsm_state198_blk = 1'b0;

    assign ap_ST_fsm_state199_blk = 1'b0;

    assign ap_ST_fsm_state19_blk  = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state200_blk = 1'b0;

    assign ap_ST_fsm_state201_blk = 1'b0;

    assign ap_ST_fsm_state202_blk = 1'b0;

    assign ap_ST_fsm_state203_blk = 1'b0;

    assign ap_ST_fsm_state204_blk = 1'b0;

    assign ap_ST_fsm_state205_blk = 1'b0;

    assign ap_ST_fsm_state206_blk = 1'b0;

    assign ap_ST_fsm_state207_blk = 1'b0;

    assign ap_ST_fsm_state208_blk = 1'b0;

    assign ap_ST_fsm_state209_blk = 1'b0;

    assign ap_ST_fsm_state20_blk  = 1'b0;

    assign ap_ST_fsm_state210_blk = 1'b0;

    assign ap_ST_fsm_state211_blk = 1'b0;

    assign ap_ST_fsm_state212_blk = 1'b0;

    assign ap_ST_fsm_state213_blk = 1'b0;

    assign ap_ST_fsm_state214_blk = 1'b0;

    assign ap_ST_fsm_state215_blk = 1'b0;

    assign ap_ST_fsm_state216_blk = 1'b0;

    assign ap_ST_fsm_state217_blk = 1'b0;

    always @(*) begin
        if ((grp_sin_or_cos_double_s_fu_421_p_done == 1'b0)) begin
            ap_ST_fsm_state218_blk = 1'b1;
        end else begin
            ap_ST_fsm_state218_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state219_blk = 1'b0;

    assign ap_ST_fsm_state21_blk  = 1'b0;

    assign ap_ST_fsm_state220_blk = 1'b0;

    assign ap_ST_fsm_state221_blk = 1'b0;

    assign ap_ST_fsm_state222_blk = 1'b0;

    assign ap_ST_fsm_state223_blk = 1'b0;

    assign ap_ST_fsm_state224_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state225_on_subcall_done)) begin
            ap_ST_fsm_state225_blk = 1'b1;
        end else begin
            ap_ST_fsm_state225_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state226_blk = 1'b0;

    always @(*) begin
        if ((grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done == 1'b0)) begin
            ap_ST_fsm_state227_blk = 1'b1;
        end else begin
            ap_ST_fsm_state227_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state228_blk = 1'b0;

    assign ap_ST_fsm_state229_blk = 1'b0;

    assign ap_ST_fsm_state22_blk  = 1'b0;

    assign ap_ST_fsm_state230_blk = 1'b0;

    assign ap_ST_fsm_state231_blk = 1'b0;

    assign ap_ST_fsm_state232_blk = 1'b0;

    assign ap_ST_fsm_state233_blk = 1'b0;

    assign ap_ST_fsm_state234_blk = 1'b0;

    assign ap_ST_fsm_state235_blk = 1'b0;

    assign ap_ST_fsm_state236_blk = 1'b0;

    assign ap_ST_fsm_state237_blk = 1'b0;

    assign ap_ST_fsm_state238_blk = 1'b0;

    assign ap_ST_fsm_state239_blk = 1'b0;

    assign ap_ST_fsm_state23_blk  = 1'b0;

    assign ap_ST_fsm_state240_blk = 1'b0;

    assign ap_ST_fsm_state241_blk = 1'b0;

    assign ap_ST_fsm_state242_blk = 1'b0;

    assign ap_ST_fsm_state243_blk = 1'b0;

    assign ap_ST_fsm_state24_blk  = 1'b0;

    assign ap_ST_fsm_state25_blk  = 1'b0;

    assign ap_ST_fsm_state26_blk  = 1'b0;

    assign ap_ST_fsm_state27_blk  = 1'b0;

    assign ap_ST_fsm_state28_blk  = 1'b0;

    assign ap_ST_fsm_state29_blk  = 1'b0;

    assign ap_ST_fsm_state2_blk   = 1'b0;

    assign ap_ST_fsm_state30_blk  = 1'b0;

    assign ap_ST_fsm_state31_blk  = 1'b0;

    assign ap_ST_fsm_state32_blk  = 1'b0;

    assign ap_ST_fsm_state33_blk  = 1'b0;

    assign ap_ST_fsm_state34_blk  = 1'b0;

    assign ap_ST_fsm_state35_blk  = 1'b0;

    assign ap_ST_fsm_state36_blk  = 1'b0;

    assign ap_ST_fsm_state37_blk  = 1'b0;

    assign ap_ST_fsm_state38_blk  = 1'b0;

    assign ap_ST_fsm_state39_blk  = 1'b0;

    assign ap_ST_fsm_state3_blk   = 1'b0;

    assign ap_ST_fsm_state40_blk  = 1'b0;

    assign ap_ST_fsm_state41_blk  = 1'b0;

    assign ap_ST_fsm_state42_blk  = 1'b0;

    assign ap_ST_fsm_state43_blk  = 1'b0;

    assign ap_ST_fsm_state44_blk  = 1'b0;

    assign ap_ST_fsm_state45_blk  = 1'b0;

    assign ap_ST_fsm_state46_blk  = 1'b0;

    assign ap_ST_fsm_state47_blk  = 1'b0;

    assign ap_ST_fsm_state48_blk  = 1'b0;

    assign ap_ST_fsm_state49_blk  = 1'b0;

    assign ap_ST_fsm_state4_blk   = 1'b0;

    assign ap_ST_fsm_state50_blk  = 1'b0;

    assign ap_ST_fsm_state51_blk  = 1'b0;

    assign ap_ST_fsm_state52_blk  = 1'b0;

    assign ap_ST_fsm_state53_blk  = 1'b0;

    assign ap_ST_fsm_state54_blk  = 1'b0;

    assign ap_ST_fsm_state55_blk  = 1'b0;

    assign ap_ST_fsm_state56_blk  = 1'b0;

    assign ap_ST_fsm_state57_blk  = 1'b0;

    assign ap_ST_fsm_state58_blk  = 1'b0;

    assign ap_ST_fsm_state59_blk  = 1'b0;

    assign ap_ST_fsm_state5_blk   = 1'b0;

    assign ap_ST_fsm_state60_blk  = 1'b0;

    assign ap_ST_fsm_state61_blk  = 1'b0;

    assign ap_ST_fsm_state62_blk  = 1'b0;

    assign ap_ST_fsm_state63_blk  = 1'b0;

    assign ap_ST_fsm_state64_blk  = 1'b0;

    assign ap_ST_fsm_state65_blk  = 1'b0;

    assign ap_ST_fsm_state66_blk  = 1'b0;

    assign ap_ST_fsm_state67_blk  = 1'b0;

    assign ap_ST_fsm_state68_blk  = 1'b0;

    assign ap_ST_fsm_state69_blk  = 1'b0;

    assign ap_ST_fsm_state6_blk   = 1'b0;

    assign ap_ST_fsm_state70_blk  = 1'b0;

    assign ap_ST_fsm_state71_blk  = 1'b0;

    assign ap_ST_fsm_state72_blk  = 1'b0;

    assign ap_ST_fsm_state73_blk  = 1'b0;

    assign ap_ST_fsm_state74_blk  = 1'b0;

    assign ap_ST_fsm_state75_blk  = 1'b0;

    assign ap_ST_fsm_state76_blk  = 1'b0;

    assign ap_ST_fsm_state77_blk  = 1'b0;

    assign ap_ST_fsm_state78_blk  = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state79_on_subcall_done)) begin
            ap_ST_fsm_state79_blk = 1'b1;
        end else begin
            ap_ST_fsm_state79_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state80_blk = 1'b0;

    assign ap_ST_fsm_state81_blk = 1'b0;

    assign ap_ST_fsm_state82_blk = 1'b0;

    assign ap_ST_fsm_state83_blk = 1'b0;

    assign ap_ST_fsm_state84_blk = 1'b0;

    assign ap_ST_fsm_state85_blk = 1'b0;

    assign ap_ST_fsm_state86_blk = 1'b0;

    assign ap_ST_fsm_state87_blk = 1'b0;

    assign ap_ST_fsm_state88_blk = 1'b0;

    assign ap_ST_fsm_state89_blk = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state90_blk = 1'b0;

    assign ap_ST_fsm_state91_blk = 1'b0;

    assign ap_ST_fsm_state92_blk = 1'b0;

    assign ap_ST_fsm_state93_blk = 1'b0;

    assign ap_ST_fsm_state94_blk = 1'b0;

    assign ap_ST_fsm_state95_blk = 1'b0;

    assign ap_ST_fsm_state96_blk = 1'b0;

    assign ap_ST_fsm_state97_blk = 1'b0;

    assign ap_ST_fsm_state98_blk = 1'b0;

    assign ap_ST_fsm_state99_blk = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if ((((1'b1 == ap_CS_fsm_state208) & ((icmp_ln134_fu_778_p2 == 1'd1) | (1'd1 == and_ln107_reg_936))) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state208) & ((icmp_ln134_fu_778_p2 == 1'd1) | (1'd1 == and_ln107_reg_936)))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_266_p0 = currOdometry_0_2_val;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_266_p0 = currOdometry_0_0_val;
        end else begin
            grp_fu_266_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_266_p1 = prevOdometry_0_2_val;
        end else if ((1'b1 == ap_CS_fsm_state1)) begin
            grp_fu_266_p1 = prevOdometry_0_0_val;
        end else begin
            grp_fu_266_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state59)) begin
            grp_fu_295_p0 = zext_ln57_1_fu_727_p1;
        end else if ((1'b1 == ap_CS_fsm_state52)) begin
            grp_fu_295_p0 = zext_ln57_4_fu_716_p1;
        end else if ((1'b1 == ap_CS_fsm_state46)) begin
            grp_fu_295_p0 = zext_ln57_2_fu_711_p1;
        end else if ((1'b1 == ap_CS_fsm_state40)) begin
            grp_fu_295_p0 = zext_ln57_fu_706_p1;
        end else begin
            grp_fu_295_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state197) | (1'b1 == ap_CS_fsm_state190))) begin
            grp_fu_304_p0 = reg_530;
        end else if ((1'b1 == ap_CS_fsm_state179)) begin
            grp_fu_304_p0 = reg_551;
        end else if ((1'b1 == ap_CS_fsm_state172)) begin
            grp_fu_304_p0 = reg_557;
        end else begin
            grp_fu_304_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state190)) begin
            grp_fu_307_p0 = reg_538;
        end else if ((1'b1 == ap_CS_fsm_state172)) begin
            grp_fu_307_p0 = scaleH2_reg_1109;
        end else begin
            grp_fu_307_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state200) | (1'b1 == ap_CS_fsm_state193) | (1'b1 == ap_CS_fsm_state182) | (1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state199) | (1'b1 == ap_CS_fsm_state192) | (1'b1 == ap_CS_fsm_state181) | (1'b1 == ap_CS_fsm_state174) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state6) | ((1'b0 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79)))) begin
            grp_fu_310_ce = 1'b1;
        end else begin
            grp_fu_310_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state199) | (1'b1 == ap_CS_fsm_state192) | (1'b1 == ap_CS_fsm_state181) | (1'b1 == ap_CS_fsm_state174))) begin
            grp_fu_310_p0 = reg_563;
        end else if ((1'b1 == ap_CS_fsm_state78)) begin
            grp_fu_310_p0 = prevOdometry_0_2_val;
        end else if (((1'b1 == ap_CS_fsm_state50) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state56))) begin
            grp_fu_310_p0 = reg_466;
        end else if (((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state6))) begin
            grp_fu_310_p0 = reg_406;
        end else begin
            grp_fu_310_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state192) | (1'b1 == ap_CS_fsm_state174))) begin
            grp_fu_313_p0 = reg_568;
        end else if ((1'b1 == ap_CS_fsm_state69)) begin
            grp_fu_313_p0 = u2_1_reg_1005;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_313_p0 = sub5_reg_889;
        end else begin
            grp_fu_313_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state217) | (1'b1 == ap_CS_fsm_state236) | (1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state210) | (1'b1 == ap_CS_fsm_state111) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state198) | (1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state223) | (1'b1 == ap_CS_fsm_state121) | (1'b1 == ap_CS_fsm_state242) | (1'b1 == ap_CS_fsm_state216) | (1'b1 == ap_CS_fsm_state196) | (1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state92) | (1'b1 == ap_CS_fsm_state207) | (1'b1 == ap_CS_fsm_state86) | (1'b1 == ap_CS_fsm_state232) | (1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state93) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state200) | (1'b1 == ap_CS_fsm_state193) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state241) | (1'b1 == ap_CS_fsm_state240) | (1'b1 == ap_CS_fsm_state239) | (1'b1 == ap_CS_fsm_state238) | (1'b1 == ap_CS_fsm_state237) | (1'b1 == ap_CS_fsm_state231) | (1'b1 == ap_CS_fsm_state230) 
    | (1'b1 == ap_CS_fsm_state229) | (1'b1 == ap_CS_fsm_state228) | (1'b1 == ap_CS_fsm_state222) | (1'b1 == ap_CS_fsm_state221) | (1'b1 == ap_CS_fsm_state220) | (1'b1 == ap_CS_fsm_state215) | (1'b1 == ap_CS_fsm_state214) | (1'b1 == ap_CS_fsm_state213) | (1'b1 == ap_CS_fsm_state212) | (1'b1 == ap_CS_fsm_state211) | (1'b1 == ap_CS_fsm_state206) | (1'b1 == ap_CS_fsm_state205) | (1'b1 == ap_CS_fsm_state204) | (1'b1 == ap_CS_fsm_state203) | (1'b1 == ap_CS_fsm_state202) | (1'b1 == ap_CS_fsm_state195) | (1'b1 == ap_CS_fsm_state188) | (1'b1 == ap_CS_fsm_state187) | (1'b1 == ap_CS_fsm_state186) | (1'b1 == ap_CS_fsm_state185) | (1'b1 == ap_CS_fsm_state184) | (1'b1 == ap_CS_fsm_state120) | (1'b1 == ap_CS_fsm_state119) | (1'b1 == ap_CS_fsm_state118) | (1'b1 == ap_CS_fsm_state117) | (1'b1 == ap_CS_fsm_state116) | (1'b1 == ap_CS_fsm_state113) | (1'b1 == ap_CS_fsm_state110) | (1'b1 == ap_CS_fsm_state109) | (1'b1 == ap_CS_fsm_state91) | (1'b1 == ap_CS_fsm_state90) | (1'b1 == ap_CS_fsm_state89) | (1'b1 == ap_CS_fsm_state88) | (1'b1 
    == ap_CS_fsm_state85) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state35) | (1'b1 == ap_CS_fsm_state34) | (1'b1 == ap_CS_fsm_state33) | (1'b1 == ap_CS_fsm_state32) | (1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state112) | (1'b1 == ap_CS_fsm_state219) | (1'b1 == ap_CS_fsm_state201) | (1'b1 == ap_CS_fsm_state194) | (1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state115) | (1'b1 == ap_CS_fsm_state108) | (1'b1 == ap_CS_fsm_state87) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state199) | (1'b1 == ap_CS_fsm_state192) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state197) | (1'b1 == ap_CS_fsm_state190) | ((grp_sin_or_cos_double_s_fu_196_ap_done 
    == 1'b1) & (1'b1 == ap_CS_fsm_state218)) | ((grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state227)))) begin
            grp_fu_319_ce = 1'b1;
        end else begin
            grp_fu_319_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state201) | (1'b1 == ap_CS_fsm_state194) | (1'b1 == ap_CS_fsm_state87) | (1'b1 == ap_CS_fsm_state80))) begin
            grp_fu_319_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state217) | (1'b1 == ap_CS_fsm_state236) | (1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state210) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state115) | (1'b1 == ap_CS_fsm_state108) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state190))) begin
            grp_fu_319_opcode = 2'd0;
        end else begin
            grp_fu_319_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state236)) begin
            grp_fu_319_p0 = bitcast_ln138_fu_826_p1;
        end else if ((1'b1 == ap_CS_fsm_state226)) begin
            grp_fu_319_p0 = bitcast_ln137_fu_809_p1;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_319_p0 = reg_530;
        end else if ((1'b1 == ap_CS_fsm_state210)) begin
            grp_fu_319_p0 = bitcast_ln135_fu_804_p1;
        end else if ((1'b1 == ap_CS_fsm_state201)) begin
            grp_fu_319_p0 = dTrans_reg_1050;
        end else if ((1'b1 == ap_CS_fsm_state194)) begin
            grp_fu_319_p0 = reg_483;
        end else if ((1'b1 == ap_CS_fsm_state115)) begin
            grp_fu_319_p0 = reg_538;
        end else if ((1'b1 == ap_CS_fsm_state108)) begin
            grp_fu_319_p0 = reg_505;
        end else if ((1'b1 == ap_CS_fsm_state87)) begin
            grp_fu_319_p0 = thetaDiff_reg_915;
        end else if ((1'b1 == ap_CS_fsm_state80)) begin
            grp_fu_319_p0 = tmp_s_reg_1030;
        end else if (((1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state190))) begin
            grp_fu_319_p0 = reg_439;
        end else if ((1'b1 == ap_CS_fsm_state15)) begin
            grp_fu_319_p0 = reg_427;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_319_p0 = bitcast_ln497_fu_610_p1;
        end else begin
            grp_fu_319_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state236) | (1'b1 == ap_CS_fsm_state226))) begin
            grp_fu_319_p1 = reg_439;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_319_p1 = reg_538;
        end else if ((1'b1 == ap_CS_fsm_state210)) begin
            grp_fu_319_p1 = reg_427;
        end else if (((1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state190))) begin
            grp_fu_319_p1 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state115)) begin
            grp_fu_319_p1 = reg_505;
        end else if ((1'b1 == ap_CS_fsm_state87)) begin
            grp_fu_319_p1 = reg_483;
        end else if (((1'b1 == ap_CS_fsm_state201) | (1'b1 == ap_CS_fsm_state194) | (1'b1 == ap_CS_fsm_state80))) begin
            grp_fu_319_p1 = reg_411;
        end else if (((1'b1 == ap_CS_fsm_state108) | (1'b1 == ap_CS_fsm_state30))) begin
            grp_fu_319_p1 = reg_448;
        end else if ((1'b1 == ap_CS_fsm_state15)) begin
            grp_fu_319_p1 = bitcast_ln497_2_fu_651_p1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            grp_fu_319_p1 = bitcast_ln497_1_fu_631_p1;
        end else begin
            grp_fu_319_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_323_ce = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_323_ce = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_323_ce = grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_ce;
        end else begin
            grp_fu_323_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_323_opcode = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_323_opcode = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_323_opcode = grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state194)) begin
            grp_fu_323_opcode = 2'd1;
        end else if (((1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state108))) begin
            grp_fu_323_opcode = 2'd0;
        end else begin
            grp_fu_323_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_323_p0 = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_323_p0 = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_323_p0 = grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state194)) begin
            grp_fu_323_p0 = reg_427;
        end else if ((1'b1 == ap_CS_fsm_state183)) begin
            grp_fu_323_p0 = reg_448;
        end else if ((1'b1 == ap_CS_fsm_state108)) begin
            grp_fu_323_p0 = reg_471;
        end else begin
            grp_fu_323_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_323_p1 = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_323_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_323_p1 = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_323_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_323_p1 = grp_atan2_cordic_double_s_fu_188_grp_fu_323_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state194)) begin
            grp_fu_323_p1 = reg_419;
        end else if ((1'b1 == ap_CS_fsm_state183)) begin
            grp_fu_323_p1 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state108)) begin
            grp_fu_323_p1 = reg_512;
        end else begin
            grp_fu_323_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state111) | (1'b1 == ap_CS_fsm_state98) | (1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state180) | (1'b1 == ap_CS_fsm_state173) | (1'b1 == ap_CS_fsm_state171) | (1'b1 == ap_CS_fsm_state162) | (1'b1 == ap_CS_fsm_state178) | (1'b1 == ap_CS_fsm_state168) | (1'b1 == ap_CS_fsm_state223) | (1'b1 == ap_CS_fsm_state105) | (1'b1 == ap_CS_fsm_state169) | (1'b1 == ap_CS_fsm_state114) | (1'b1 == ap_CS_fsm_state104) | (1'b1 == ap_CS_fsm_state107) | (1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state232) | (1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state163) | (1'b1 == ap_CS_fsm_state99) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state93) | (1'b1 == ap_CS_fsm_state182) | (1'b1 == ap_CS_fsm_state175) | (1'b1 == ap_CS_fsm_state177) | (1'b1 == ap_CS_fsm_state170) | (1'b1 == ap_CS_fsm_state167) | (1'b1 == ap_CS_fsm_state166) | (1'b1 == ap_CS_fsm_state165) | (1'b1 == ap_CS_fsm_state164) | (1'b1 == 
    ap_CS_fsm_state161) | (1'b1 == ap_CS_fsm_state160) | (1'b1 == ap_CS_fsm_state159) | (1'b1 == ap_CS_fsm_state158) | (1'b1 == ap_CS_fsm_state103) | (1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state97) | (1'b1 == ap_CS_fsm_state96) | (1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state76) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state231) | (1'b1 == ap_CS_fsm_state230) | (1'b1 == ap_CS_fsm_state229) | (1'b1 == ap_CS_fsm_state228) | (1'b1 == ap_CS_fsm_state222) | (1'b1 == ap_CS_fsm_state221) | (1'b1 == ap_CS_fsm_state220) | (1'b1 == ap_CS_fsm_state188) | (1'b1 == ap_CS_fsm_state187) | (1'b1 == ap_CS_fsm_state186) | (1'b1 == ap_CS_fsm_state185) | (1'b1 == ap_CS_fsm_state184) | (1'b1 == ap_CS_fsm_state113) | (1'b1 == ap_CS_fsm_state110) | (1'b1 == ap_CS_fsm_state109) | (1'b1 == ap_CS_fsm_state112) 
    | (1'b1 == ap_CS_fsm_state106) | (1'b1 == ap_CS_fsm_state219) | (1'b1 == ap_CS_fsm_state176) | (1'b1 == ap_CS_fsm_state157) | (1'b1 == ap_CS_fsm_state101) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state108) | (1'b1 == ap_CS_fsm_state181) | (1'b1 == ap_CS_fsm_state174) | (1'b1 == ap_CS_fsm_state179) | (1'b1 == ap_CS_fsm_state172) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state224) | ((1'b0 == ap_block_state225_on_subcall_done) & (1'b1 == ap_CS_fsm_state225)) | ((grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state227)))) begin
            grp_fu_333_ce = 1'b1;
        end else begin
            grp_fu_333_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state219))) begin
            grp_fu_333_p0 = reg_483;
        end else if ((1'b1 == ap_CS_fsm_state176)) begin
            grp_fu_333_p0 = reg_439;
        end else if ((1'b1 == ap_CS_fsm_state163)) begin
            grp_fu_333_p0 = reg_557;
        end else if (((1'b1 == ap_CS_fsm_state169) | (1'b1 == ap_CS_fsm_state157))) begin
            grp_fu_333_p0 = reg_551;
        end else if ((1'b1 == ap_CS_fsm_state108)) begin
            grp_fu_333_p0 = reg_518;
        end else if (((1'b1 == ap_CS_fsm_state101) | (1'b1 == ap_CS_fsm_state183))) begin
            grp_fu_333_p0 = reg_505;
        end else if ((1'b1 == ap_CS_fsm_state99)) begin
            grp_fu_333_p0 = tmp_16_reg_1089;
        end else if ((1'b1 == ap_CS_fsm_state94)) begin
            grp_fu_333_p0 = bitcast_ln116_fu_756_p1;
        end else if (((1'b1 == ap_CS_fsm_state105) | (1'b1 == ap_CS_fsm_state93))) begin
            grp_fu_333_p0 = reg_492;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_333_p0 = conv3_i_reg_1015;
        end else if ((1'b1 == ap_CS_fsm_state23)) begin
            grp_fu_333_p0 = reg_411;
        end else begin
            grp_fu_333_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state169)) begin
            grp_fu_333_p1 = tmp_21_reg_1040;
        end else if ((1'b1 == ap_CS_fsm_state163)) begin
            grp_fu_333_p1 = tmp_18_reg_1035;
        end else if (((1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state219) | (1'b1 == ap_CS_fsm_state157))) begin
            grp_fu_333_p1 = reg_478;
        end else if ((1'b1 == ap_CS_fsm_state108)) begin
            grp_fu_333_p1 = reg_427;
        end else if (((1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state101))) begin
            grp_fu_333_p1 = reg_483;
        end else if (((1'b1 == ap_CS_fsm_state105) | (1'b1 == ap_CS_fsm_state99) | (1'b1 == ap_CS_fsm_state93))) begin
            grp_fu_333_p1 = 64'd13835058055282163712;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_333_p1 = 64'd4618760256179416344;
        end else if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state176) | (1'b1 == ap_CS_fsm_state183))) begin
            grp_fu_333_p1 = reg_411;
        end else begin
            grp_fu_333_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state176)) begin
            grp_fu_337_p0 = reg_524;
        end else if ((1'b1 == ap_CS_fsm_state101)) begin
            grp_fu_337_p0 = reg_448;
        end else if ((1'b1 == ap_CS_fsm_state94)) begin
            grp_fu_337_p0 = bitcast_ln116_1_fu_761_p1;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_337_p0 = conv3_i1_reg_1020;
        end else if ((1'b1 == ap_CS_fsm_state23)) begin
            grp_fu_337_p0 = reg_419;
        end else begin
            grp_fu_337_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state101))) begin
            grp_fu_337_p1 = dTrans_reg_1050;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_337_p1 = 64'd4618760256179416344;
        end else if (((1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state176))) begin
            grp_fu_337_p1 = reg_419;
        end else begin
            grp_fu_337_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state101)) begin
            grp_fu_343_p0 = reg_471;
        end else if ((1'b1 == ap_CS_fsm_state94)) begin
            grp_fu_343_p0 = bitcast_ln117_fu_766_p1;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_343_p0 = conv3_i2_reg_1025;
        end else begin
            grp_fu_343_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state101))) begin
            grp_fu_343_p1 = dTrans_reg_1050;
        end else if ((1'b1 == ap_CS_fsm_state71)) begin
            grp_fu_343_p1 = 64'd4618760256179416344;
        end else begin
            grp_fu_343_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state101)) begin
            grp_fu_349_p0 = reg_512;
        end else if ((1'b1 == ap_CS_fsm_state94)) begin
            grp_fu_349_p0 = bitcast_ln117_1_fu_771_p1;
        end else begin
            grp_fu_349_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state101)) begin
            grp_fu_353_p0 = bitcast_ln117_1_reg_1083;
        end else if ((1'b1 == ap_CS_fsm_state94)) begin
            grp_fu_353_p0 = bitcast_ln116_fu_756_p1;
        end else begin
            grp_fu_353_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_361_ce = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_361_ce = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_361_ce = grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_ce;
        end else begin
            grp_fu_361_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_361_opcode = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_361_opcode = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_361_opcode = grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_361_opcode = 5'd4;
        end else begin
            grp_fu_361_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_361_p0 = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_361_p0 = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_361_p0 = grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_361_p0 = reg_427;
        end else begin
            grp_fu_361_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state227)) begin
            grp_fu_361_p1 = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_grp_fu_361_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_fu_361_p1 = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_grp_fu_361_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_fu_361_p1 = grp_atan2_cordic_double_s_fu_188_grp_fu_361_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_361_p1 = 64'd4457293557087583675;
        end else begin
            grp_fu_361_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state217) | (1'b1 == ap_CS_fsm_state236) | (1'b1 == ap_CS_fsm_state226) | (1'b1 == ap_CS_fsm_state210) | (1'b1 == ap_CS_fsm_state208) | (1'b1 == ap_CS_fsm_state98) | (1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state198) | (1'b1 == ap_CS_fsm_state191) | (1'b1 == ap_CS_fsm_state180) | (1'b1 == ap_CS_fsm_state223) | (1'b1 == ap_CS_fsm_state242) | (1'b1 == ap_CS_fsm_state216) | (1'b1 == ap_CS_fsm_state196) | (1'b1 == ap_CS_fsm_state209) | (1'b1 == ap_CS_fsm_state235) | (1'b1 == ap_CS_fsm_state207) | (1'b1 == ap_CS_fsm_state218) | (1'b1 == ap_CS_fsm_state232) | (1'b1 == ap_CS_fsm_state225) | (1'b1 == ap_CS_fsm_state189) | (1'b1 == ap_CS_fsm_state99) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state200) | (1'b1 == ap_CS_fsm_state193) | (1'b1 == ap_CS_fsm_state182) | (1'b1 == ap_CS_fsm_state7) 
    | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state1) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state97) | (1'b1 == ap_CS_fsm_state96) | (1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state241) | (1'b1 == ap_CS_fsm_state240) | (1'b1 == ap_CS_fsm_state239) | (1'b1 == ap_CS_fsm_state238) | (1'b1 == ap_CS_fsm_state237) | (1'b1 == ap_CS_fsm_state231) | (1'b1 == ap_CS_fsm_state230) | (1'b1 == ap_CS_fsm_state229) | (1'b1 == ap_CS_fsm_state228) | (1'b1 == ap_CS_fsm_state222) | (1'b1 == ap_CS_fsm_state221) | (1'b1 == ap_CS_fsm_state220) | (1'b1 == ap_CS_fsm_state215) | (1'b1 == ap_CS_fsm_state214) | (1'b1 == ap_CS_fsm_state213) | (1'b1 == ap_CS_fsm_state212) | (1'b1 == ap_CS_fsm_state211) | (1'b1 == ap_CS_fsm_state206) | (1'b1 == ap_CS_fsm_state205) | (1'b1 == ap_CS_fsm_state204) | (1'b1 == ap_CS_fsm_state203) 
    | (1'b1 == ap_CS_fsm_state202) | (1'b1 == ap_CS_fsm_state195) | (1'b1 == ap_CS_fsm_state188) | (1'b1 == ap_CS_fsm_state187) | (1'b1 == ap_CS_fsm_state186) | (1'b1 == ap_CS_fsm_state185) | (1'b1 == ap_CS_fsm_state184) | (1'b1 == ap_CS_fsm_state35) | (1'b1 == ap_CS_fsm_state34) | (1'b1 == ap_CS_fsm_state33) | (1'b1 == ap_CS_fsm_state32) | (1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state219) | (1'b1 == ap_CS_fsm_state201) | (1'b1 == ap_CS_fsm_state194) | (1'b1 == ap_CS_fsm_state183) | (1'b1 == ap_CS_fsm_state30) | (1'b1 == ap_CS_fsm_state199) | (1'b1 == ap_CS_fsm_state192) | (1'b1 == ap_CS_fsm_state181) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state197) | (1'b1 == ap_CS_fsm_state190) | (1'b1 == ap_CS_fsm_state179) | (1'b1 == ap_CS_fsm_state234) 
    | (1'b1 == ap_CS_fsm_state233) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state243) | (1'b1 == ap_CS_fsm_state227) | (1'b1 == ap_CS_fsm_state224) | ((1'b1 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79)))) begin
            grp_fu_366_ce = 1'b0;
        end else begin
            grp_fu_366_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state122)) begin
            grp_fu_366_p1 = reg_545;
        end else if ((1'b1 == ap_CS_fsm_state115)) begin
            grp_fu_366_p1 = reg_530;
        end else if ((1'b1 == ap_CS_fsm_state112)) begin
            grp_fu_366_p1 = mul_i2_reg_1099;
        end else if ((1'b1 == ap_CS_fsm_state106)) begin
            grp_fu_366_p1 = reg_524;
        end else if ((1'b1 == ap_CS_fsm_state100)) begin
            grp_fu_366_p1 = reg_439;
        end else if ((1'b1 == ap_CS_fsm_state37)) begin
            grp_fu_366_p1 = reg_427;
        end else begin
            grp_fu_366_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state98) | (1'b1 == ap_CS_fsm_state94) | (1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state58) | (1'b1 == ap_CS_fsm_state104) | (1'b1 == ap_CS_fsm_state92) | (1'b1 == ap_CS_fsm_state86) | (1'b1 == ap_CS_fsm_state68) | (1'b1 == ap_CS_fsm_state61) | (1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state99) | (1'b1 == ap_CS_fsm_state77) | (1'b1 == ap_CS_fsm_state93) | (1'b1 == ap_CS_fsm_state67) | (1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state54) | (1'b1 == ap_CS_fsm_state53) | (1'b1 == ap_CS_fsm_state103) | (1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state97) | (1'b1 == ap_CS_fsm_state96) | (1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state76) | (1'b1 == ap_CS_fsm_state75) | (1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73) | 
    (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state91) | (1'b1 == ap_CS_fsm_state90) | (1'b1 == ap_CS_fsm_state89) | (1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state85) | (1'b1 == ap_CS_fsm_state84) | (1'b1 == ap_CS_fsm_state83) | (1'b1 == ap_CS_fsm_state82) | (1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state101) | (1'b1 == ap_CS_fsm_state71) | (1'b1 == ap_CS_fsm_state87) | (1'b1 == ap_CS_fsm_state80) | (1'b1 == ap_CS_fsm_state69) | (1'b1 == ap_CS_fsm_state62) | (1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state65) | ((1'b0 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79)))) begin
            grp_fu_376_ce = 1'b1;
        end else begin
            grp_fu_376_ce = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state64)) begin
            grp_fu_376_p1 = conv2_i2_reg_990;
        end else if ((1'b1 == ap_CS_fsm_state58)) begin
            grp_fu_376_p1 = conv2_i1_reg_970;
        end else if ((1'b1 == ap_CS_fsm_state52)) begin
            grp_fu_376_p1 = conv2_i_reg_960;
        end else begin
            grp_fu_376_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state56)) begin
            grp_fu_381_p0 = reg_589;
        end else if (((1'b1 == ap_CS_fsm_state46) | (1'b1 == ap_CS_fsm_state49))) begin
            grp_fu_381_p0 = reg_584;
        end else if (((1'b1 == ap_CS_fsm_state40) | (1'b1 == ap_CS_fsm_state43))) begin
            grp_fu_381_p0 = reg_579;
        end else if ((1'b1 == ap_CS_fsm_state37)) begin
            grp_fu_381_p0 = seed;
        end else begin
            grp_fu_381_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state225)) begin
            grp_sin_or_cos_double_s_fu_196_do_cos = 1'd0;
        end else if (((1'b1 == ap_CS_fsm_state218) | (1'b1 == ap_CS_fsm_state79))) begin
            grp_sin_or_cos_double_s_fu_196_do_cos = 1'd1;
        end else begin
            grp_sin_or_cos_double_s_fu_196_do_cos = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state218) | (1'b1 == ap_CS_fsm_state225))) begin
            grp_sin_or_cos_double_s_fu_196_t_in = reg_530;
        end else if ((1'b1 == ap_CS_fsm_state79)) begin
            grp_sin_or_cos_double_s_fu_196_t_in = reg_439;
        end else begin
            grp_sin_or_cos_double_s_fu_196_t_in = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state234) | (1'b1 == ap_CS_fsm_state233) | (1'b1 == ap_CS_fsm_state243))) begin
            pf_address0 = pf_addr_4_reg_1117;
        end else if ((1'b1 == ap_CS_fsm_state208)) begin
            pf_address0 = zext_ln134_fu_790_p1;
        end else if ((1'b1 == ap_CS_fsm_state92)) begin
            pf_address0 = 64'd80500;
        end else begin
            pf_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state208) | (1'b1 == ap_CS_fsm_state92) | (1'b1 == ap_CS_fsm_state234) | (1'b1 == ap_CS_fsm_state233) | (1'b1 == ap_CS_fsm_state243))) begin
            pf_ce0 = 1'b1;
        end else begin
            pf_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state243)) begin
            pf_d0 = zext_ln139_fu_852_p1;
        end else if ((1'b1 == ap_CS_fsm_state233)) begin
            pf_d0 = zext_ln137_fu_821_p1;
        end else begin
            pf_d0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state243)) begin
            pf_we0 = 32'd16776960;
        end else if ((1'b1 == ap_CS_fsm_state233)) begin
            pf_we0 = 32'd255;
        end else begin
            pf_we0 = 32'd0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                if (((1'b1 == ap_CS_fsm_state23) & (1'd1 == and_ln107_fu_690_p2))) begin
                    ap_NS_fsm = ap_ST_fsm_state208;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state24;
                end
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end
            ap_ST_fsm_state78: begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
            ap_ST_fsm_state79: begin
                if (((1'b0 == ap_block_state79_on_subcall_done) & (1'b1 == ap_CS_fsm_state79))) begin
                    ap_NS_fsm = ap_ST_fsm_state80;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state79;
                end
            end
            ap_ST_fsm_state80: begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
            ap_ST_fsm_state81: begin
                ap_NS_fsm = ap_ST_fsm_state82;
            end
            ap_ST_fsm_state82: begin
                ap_NS_fsm = ap_ST_fsm_state83;
            end
            ap_ST_fsm_state83: begin
                ap_NS_fsm = ap_ST_fsm_state84;
            end
            ap_ST_fsm_state84: begin
                ap_NS_fsm = ap_ST_fsm_state85;
            end
            ap_ST_fsm_state85: begin
                ap_NS_fsm = ap_ST_fsm_state86;
            end
            ap_ST_fsm_state86: begin
                ap_NS_fsm = ap_ST_fsm_state87;
            end
            ap_ST_fsm_state87: begin
                ap_NS_fsm = ap_ST_fsm_state88;
            end
            ap_ST_fsm_state88: begin
                ap_NS_fsm = ap_ST_fsm_state89;
            end
            ap_ST_fsm_state89: begin
                ap_NS_fsm = ap_ST_fsm_state90;
            end
            ap_ST_fsm_state90: begin
                ap_NS_fsm = ap_ST_fsm_state91;
            end
            ap_ST_fsm_state91: begin
                ap_NS_fsm = ap_ST_fsm_state92;
            end
            ap_ST_fsm_state92: begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end
            ap_ST_fsm_state93: begin
                ap_NS_fsm = ap_ST_fsm_state94;
            end
            ap_ST_fsm_state94: begin
                ap_NS_fsm = ap_ST_fsm_state95;
            end
            ap_ST_fsm_state95: begin
                ap_NS_fsm = ap_ST_fsm_state96;
            end
            ap_ST_fsm_state96: begin
                ap_NS_fsm = ap_ST_fsm_state97;
            end
            ap_ST_fsm_state97: begin
                ap_NS_fsm = ap_ST_fsm_state98;
            end
            ap_ST_fsm_state98: begin
                ap_NS_fsm = ap_ST_fsm_state99;
            end
            ap_ST_fsm_state99: begin
                ap_NS_fsm = ap_ST_fsm_state100;
            end
            ap_ST_fsm_state100: begin
                ap_NS_fsm = ap_ST_fsm_state101;
            end
            ap_ST_fsm_state101: begin
                ap_NS_fsm = ap_ST_fsm_state102;
            end
            ap_ST_fsm_state102: begin
                ap_NS_fsm = ap_ST_fsm_state103;
            end
            ap_ST_fsm_state103: begin
                ap_NS_fsm = ap_ST_fsm_state104;
            end
            ap_ST_fsm_state104: begin
                ap_NS_fsm = ap_ST_fsm_state105;
            end
            ap_ST_fsm_state105: begin
                ap_NS_fsm = ap_ST_fsm_state106;
            end
            ap_ST_fsm_state106: begin
                ap_NS_fsm = ap_ST_fsm_state107;
            end
            ap_ST_fsm_state107: begin
                ap_NS_fsm = ap_ST_fsm_state108;
            end
            ap_ST_fsm_state108: begin
                ap_NS_fsm = ap_ST_fsm_state109;
            end
            ap_ST_fsm_state109: begin
                ap_NS_fsm = ap_ST_fsm_state110;
            end
            ap_ST_fsm_state110: begin
                ap_NS_fsm = ap_ST_fsm_state111;
            end
            ap_ST_fsm_state111: begin
                ap_NS_fsm = ap_ST_fsm_state112;
            end
            ap_ST_fsm_state112: begin
                ap_NS_fsm = ap_ST_fsm_state113;
            end
            ap_ST_fsm_state113: begin
                ap_NS_fsm = ap_ST_fsm_state114;
            end
            ap_ST_fsm_state114: begin
                ap_NS_fsm = ap_ST_fsm_state115;
            end
            ap_ST_fsm_state115: begin
                ap_NS_fsm = ap_ST_fsm_state116;
            end
            ap_ST_fsm_state116: begin
                ap_NS_fsm = ap_ST_fsm_state117;
            end
            ap_ST_fsm_state117: begin
                ap_NS_fsm = ap_ST_fsm_state118;
            end
            ap_ST_fsm_state118: begin
                ap_NS_fsm = ap_ST_fsm_state119;
            end
            ap_ST_fsm_state119: begin
                ap_NS_fsm = ap_ST_fsm_state120;
            end
            ap_ST_fsm_state120: begin
                ap_NS_fsm = ap_ST_fsm_state121;
            end
            ap_ST_fsm_state121: begin
                ap_NS_fsm = ap_ST_fsm_state122;
            end
            ap_ST_fsm_state122: begin
                ap_NS_fsm = ap_ST_fsm_state123;
            end
            ap_ST_fsm_state123: begin
                ap_NS_fsm = ap_ST_fsm_state124;
            end
            ap_ST_fsm_state124: begin
                ap_NS_fsm = ap_ST_fsm_state125;
            end
            ap_ST_fsm_state125: begin
                ap_NS_fsm = ap_ST_fsm_state126;
            end
            ap_ST_fsm_state126: begin
                ap_NS_fsm = ap_ST_fsm_state127;
            end
            ap_ST_fsm_state127: begin
                ap_NS_fsm = ap_ST_fsm_state128;
            end
            ap_ST_fsm_state128: begin
                ap_NS_fsm = ap_ST_fsm_state129;
            end
            ap_ST_fsm_state129: begin
                ap_NS_fsm = ap_ST_fsm_state130;
            end
            ap_ST_fsm_state130: begin
                ap_NS_fsm = ap_ST_fsm_state131;
            end
            ap_ST_fsm_state131: begin
                ap_NS_fsm = ap_ST_fsm_state132;
            end
            ap_ST_fsm_state132: begin
                ap_NS_fsm = ap_ST_fsm_state133;
            end
            ap_ST_fsm_state133: begin
                ap_NS_fsm = ap_ST_fsm_state134;
            end
            ap_ST_fsm_state134: begin
                ap_NS_fsm = ap_ST_fsm_state135;
            end
            ap_ST_fsm_state135: begin
                ap_NS_fsm = ap_ST_fsm_state136;
            end
            ap_ST_fsm_state136: begin
                ap_NS_fsm = ap_ST_fsm_state137;
            end
            ap_ST_fsm_state137: begin
                ap_NS_fsm = ap_ST_fsm_state138;
            end
            ap_ST_fsm_state138: begin
                ap_NS_fsm = ap_ST_fsm_state139;
            end
            ap_ST_fsm_state139: begin
                ap_NS_fsm = ap_ST_fsm_state140;
            end
            ap_ST_fsm_state140: begin
                ap_NS_fsm = ap_ST_fsm_state141;
            end
            ap_ST_fsm_state141: begin
                ap_NS_fsm = ap_ST_fsm_state142;
            end
            ap_ST_fsm_state142: begin
                ap_NS_fsm = ap_ST_fsm_state143;
            end
            ap_ST_fsm_state143: begin
                ap_NS_fsm = ap_ST_fsm_state144;
            end
            ap_ST_fsm_state144: begin
                ap_NS_fsm = ap_ST_fsm_state145;
            end
            ap_ST_fsm_state145: begin
                ap_NS_fsm = ap_ST_fsm_state146;
            end
            ap_ST_fsm_state146: begin
                ap_NS_fsm = ap_ST_fsm_state147;
            end
            ap_ST_fsm_state147: begin
                ap_NS_fsm = ap_ST_fsm_state148;
            end
            ap_ST_fsm_state148: begin
                ap_NS_fsm = ap_ST_fsm_state149;
            end
            ap_ST_fsm_state149: begin
                ap_NS_fsm = ap_ST_fsm_state150;
            end
            ap_ST_fsm_state150: begin
                ap_NS_fsm = ap_ST_fsm_state151;
            end
            ap_ST_fsm_state151: begin
                ap_NS_fsm = ap_ST_fsm_state152;
            end
            ap_ST_fsm_state152: begin
                ap_NS_fsm = ap_ST_fsm_state153;
            end
            ap_ST_fsm_state153: begin
                ap_NS_fsm = ap_ST_fsm_state154;
            end
            ap_ST_fsm_state154: begin
                ap_NS_fsm = ap_ST_fsm_state155;
            end
            ap_ST_fsm_state155: begin
                ap_NS_fsm = ap_ST_fsm_state156;
            end
            ap_ST_fsm_state156: begin
                ap_NS_fsm = ap_ST_fsm_state157;
            end
            ap_ST_fsm_state157: begin
                ap_NS_fsm = ap_ST_fsm_state158;
            end
            ap_ST_fsm_state158: begin
                ap_NS_fsm = ap_ST_fsm_state159;
            end
            ap_ST_fsm_state159: begin
                ap_NS_fsm = ap_ST_fsm_state160;
            end
            ap_ST_fsm_state160: begin
                ap_NS_fsm = ap_ST_fsm_state161;
            end
            ap_ST_fsm_state161: begin
                ap_NS_fsm = ap_ST_fsm_state162;
            end
            ap_ST_fsm_state162: begin
                ap_NS_fsm = ap_ST_fsm_state163;
            end
            ap_ST_fsm_state163: begin
                ap_NS_fsm = ap_ST_fsm_state164;
            end
            ap_ST_fsm_state164: begin
                ap_NS_fsm = ap_ST_fsm_state165;
            end
            ap_ST_fsm_state165: begin
                ap_NS_fsm = ap_ST_fsm_state166;
            end
            ap_ST_fsm_state166: begin
                ap_NS_fsm = ap_ST_fsm_state167;
            end
            ap_ST_fsm_state167: begin
                ap_NS_fsm = ap_ST_fsm_state168;
            end
            ap_ST_fsm_state168: begin
                ap_NS_fsm = ap_ST_fsm_state169;
            end
            ap_ST_fsm_state169: begin
                ap_NS_fsm = ap_ST_fsm_state170;
            end
            ap_ST_fsm_state170: begin
                ap_NS_fsm = ap_ST_fsm_state171;
            end
            ap_ST_fsm_state171: begin
                ap_NS_fsm = ap_ST_fsm_state172;
            end
            ap_ST_fsm_state172: begin
                ap_NS_fsm = ap_ST_fsm_state173;
            end
            ap_ST_fsm_state173: begin
                ap_NS_fsm = ap_ST_fsm_state174;
            end
            ap_ST_fsm_state174: begin
                ap_NS_fsm = ap_ST_fsm_state175;
            end
            ap_ST_fsm_state175: begin
                ap_NS_fsm = ap_ST_fsm_state176;
            end
            ap_ST_fsm_state176: begin
                ap_NS_fsm = ap_ST_fsm_state177;
            end
            ap_ST_fsm_state177: begin
                ap_NS_fsm = ap_ST_fsm_state178;
            end
            ap_ST_fsm_state178: begin
                ap_NS_fsm = ap_ST_fsm_state179;
            end
            ap_ST_fsm_state179: begin
                ap_NS_fsm = ap_ST_fsm_state180;
            end
            ap_ST_fsm_state180: begin
                ap_NS_fsm = ap_ST_fsm_state181;
            end
            ap_ST_fsm_state181: begin
                ap_NS_fsm = ap_ST_fsm_state182;
            end
            ap_ST_fsm_state182: begin
                ap_NS_fsm = ap_ST_fsm_state183;
            end
            ap_ST_fsm_state183: begin
                ap_NS_fsm = ap_ST_fsm_state184;
            end
            ap_ST_fsm_state184: begin
                ap_NS_fsm = ap_ST_fsm_state185;
            end
            ap_ST_fsm_state185: begin
                ap_NS_fsm = ap_ST_fsm_state186;
            end
            ap_ST_fsm_state186: begin
                ap_NS_fsm = ap_ST_fsm_state187;
            end
            ap_ST_fsm_state187: begin
                ap_NS_fsm = ap_ST_fsm_state188;
            end
            ap_ST_fsm_state188: begin
                ap_NS_fsm = ap_ST_fsm_state189;
            end
            ap_ST_fsm_state189: begin
                ap_NS_fsm = ap_ST_fsm_state190;
            end
            ap_ST_fsm_state190: begin
                ap_NS_fsm = ap_ST_fsm_state191;
            end
            ap_ST_fsm_state191: begin
                ap_NS_fsm = ap_ST_fsm_state192;
            end
            ap_ST_fsm_state192: begin
                ap_NS_fsm = ap_ST_fsm_state193;
            end
            ap_ST_fsm_state193: begin
                ap_NS_fsm = ap_ST_fsm_state194;
            end
            ap_ST_fsm_state194: begin
                ap_NS_fsm = ap_ST_fsm_state195;
            end
            ap_ST_fsm_state195: begin
                ap_NS_fsm = ap_ST_fsm_state196;
            end
            ap_ST_fsm_state196: begin
                ap_NS_fsm = ap_ST_fsm_state197;
            end
            ap_ST_fsm_state197: begin
                ap_NS_fsm = ap_ST_fsm_state198;
            end
            ap_ST_fsm_state198: begin
                ap_NS_fsm = ap_ST_fsm_state199;
            end
            ap_ST_fsm_state199: begin
                ap_NS_fsm = ap_ST_fsm_state200;
            end
            ap_ST_fsm_state200: begin
                ap_NS_fsm = ap_ST_fsm_state201;
            end
            ap_ST_fsm_state201: begin
                ap_NS_fsm = ap_ST_fsm_state202;
            end
            ap_ST_fsm_state202: begin
                ap_NS_fsm = ap_ST_fsm_state203;
            end
            ap_ST_fsm_state203: begin
                ap_NS_fsm = ap_ST_fsm_state204;
            end
            ap_ST_fsm_state204: begin
                ap_NS_fsm = ap_ST_fsm_state205;
            end
            ap_ST_fsm_state205: begin
                ap_NS_fsm = ap_ST_fsm_state206;
            end
            ap_ST_fsm_state206: begin
                ap_NS_fsm = ap_ST_fsm_state207;
            end
            ap_ST_fsm_state207: begin
                ap_NS_fsm = ap_ST_fsm_state208;
            end
            ap_ST_fsm_state208: begin
                if (((1'b1 == ap_CS_fsm_state208) & ((icmp_ln134_fu_778_p2 == 1'd1) | (1'd1 == and_ln107_reg_936)))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state209;
                end
            end
            ap_ST_fsm_state209: begin
                ap_NS_fsm = ap_ST_fsm_state210;
            end
            ap_ST_fsm_state210: begin
                ap_NS_fsm = ap_ST_fsm_state211;
            end
            ap_ST_fsm_state211: begin
                ap_NS_fsm = ap_ST_fsm_state212;
            end
            ap_ST_fsm_state212: begin
                ap_NS_fsm = ap_ST_fsm_state213;
            end
            ap_ST_fsm_state213: begin
                ap_NS_fsm = ap_ST_fsm_state214;
            end
            ap_ST_fsm_state214: begin
                ap_NS_fsm = ap_ST_fsm_state215;
            end
            ap_ST_fsm_state215: begin
                ap_NS_fsm = ap_ST_fsm_state216;
            end
            ap_ST_fsm_state216: begin
                ap_NS_fsm = ap_ST_fsm_state217;
            end
            ap_ST_fsm_state217: begin
                ap_NS_fsm = ap_ST_fsm_state218;
            end
            ap_ST_fsm_state218: begin
                if (((grp_sin_or_cos_double_s_fu_196_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state218))) begin
                    ap_NS_fsm = ap_ST_fsm_state219;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state218;
                end
            end
            ap_ST_fsm_state219: begin
                ap_NS_fsm = ap_ST_fsm_state220;
            end
            ap_ST_fsm_state220: begin
                ap_NS_fsm = ap_ST_fsm_state221;
            end
            ap_ST_fsm_state221: begin
                ap_NS_fsm = ap_ST_fsm_state222;
            end
            ap_ST_fsm_state222: begin
                ap_NS_fsm = ap_ST_fsm_state223;
            end
            ap_ST_fsm_state223: begin
                ap_NS_fsm = ap_ST_fsm_state224;
            end
            ap_ST_fsm_state224: begin
                ap_NS_fsm = ap_ST_fsm_state225;
            end
            ap_ST_fsm_state225: begin
                if (((1'b0 == ap_block_state225_on_subcall_done) & (1'b1 == ap_CS_fsm_state225))) begin
                    ap_NS_fsm = ap_ST_fsm_state226;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state225;
                end
            end
            ap_ST_fsm_state226: begin
                ap_NS_fsm = ap_ST_fsm_state227;
            end
            ap_ST_fsm_state227: begin
                if (((grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state227))) begin
                    ap_NS_fsm = ap_ST_fsm_state228;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state227;
                end
            end
            ap_ST_fsm_state228: begin
                ap_NS_fsm = ap_ST_fsm_state229;
            end
            ap_ST_fsm_state229: begin
                ap_NS_fsm = ap_ST_fsm_state230;
            end
            ap_ST_fsm_state230: begin
                ap_NS_fsm = ap_ST_fsm_state231;
            end
            ap_ST_fsm_state231: begin
                ap_NS_fsm = ap_ST_fsm_state232;
            end
            ap_ST_fsm_state232: begin
                ap_NS_fsm = ap_ST_fsm_state233;
            end
            ap_ST_fsm_state233: begin
                ap_NS_fsm = ap_ST_fsm_state234;
            end
            ap_ST_fsm_state234: begin
                ap_NS_fsm = ap_ST_fsm_state235;
            end
            ap_ST_fsm_state235: begin
                ap_NS_fsm = ap_ST_fsm_state236;
            end
            ap_ST_fsm_state236: begin
                ap_NS_fsm = ap_ST_fsm_state237;
            end
            ap_ST_fsm_state237: begin
                ap_NS_fsm = ap_ST_fsm_state238;
            end
            ap_ST_fsm_state238: begin
                ap_NS_fsm = ap_ST_fsm_state239;
            end
            ap_ST_fsm_state239: begin
                ap_NS_fsm = ap_ST_fsm_state240;
            end
            ap_ST_fsm_state240: begin
                ap_NS_fsm = ap_ST_fsm_state241;
            end
            ap_ST_fsm_state241: begin
                ap_NS_fsm = ap_ST_fsm_state242;
            end
            ap_ST_fsm_state242: begin
                ap_NS_fsm = ap_ST_fsm_state243;
            end
            ap_ST_fsm_state243: begin
                ap_NS_fsm = ap_ST_fsm_state208;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln134_fu_784_p2 = (i_fu_126 + 9'd1);

    assign and_ln107_fu_690_p2 = (or_ln107_fu_686_p2 & grp_fu_413_p_dout0);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state100 = ap_CS_fsm[32'd99];

    assign ap_CS_fsm_state101 = ap_CS_fsm[32'd100];

    assign ap_CS_fsm_state102 = ap_CS_fsm[32'd101];

    assign ap_CS_fsm_state103 = ap_CS_fsm[32'd102];

    assign ap_CS_fsm_state104 = ap_CS_fsm[32'd103];

    assign ap_CS_fsm_state105 = ap_CS_fsm[32'd104];

    assign ap_CS_fsm_state106 = ap_CS_fsm[32'd105];

    assign ap_CS_fsm_state107 = ap_CS_fsm[32'd106];

    assign ap_CS_fsm_state108 = ap_CS_fsm[32'd107];

    assign ap_CS_fsm_state109 = ap_CS_fsm[32'd108];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state110 = ap_CS_fsm[32'd109];

    assign ap_CS_fsm_state111 = ap_CS_fsm[32'd110];

    assign ap_CS_fsm_state112 = ap_CS_fsm[32'd111];

    assign ap_CS_fsm_state113 = ap_CS_fsm[32'd112];

    assign ap_CS_fsm_state114 = ap_CS_fsm[32'd113];

    assign ap_CS_fsm_state115 = ap_CS_fsm[32'd114];

    assign ap_CS_fsm_state116 = ap_CS_fsm[32'd115];

    assign ap_CS_fsm_state117 = ap_CS_fsm[32'd116];

    assign ap_CS_fsm_state118 = ap_CS_fsm[32'd117];

    assign ap_CS_fsm_state119 = ap_CS_fsm[32'd118];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state120 = ap_CS_fsm[32'd119];

    assign ap_CS_fsm_state121 = ap_CS_fsm[32'd120];

    assign ap_CS_fsm_state122 = ap_CS_fsm[32'd121];

    assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state156 = ap_CS_fsm[32'd155];

    assign ap_CS_fsm_state157 = ap_CS_fsm[32'd156];

    assign ap_CS_fsm_state158 = ap_CS_fsm[32'd157];

    assign ap_CS_fsm_state159 = ap_CS_fsm[32'd158];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state160 = ap_CS_fsm[32'd159];

    assign ap_CS_fsm_state161 = ap_CS_fsm[32'd160];

    assign ap_CS_fsm_state162 = ap_CS_fsm[32'd161];

    assign ap_CS_fsm_state163 = ap_CS_fsm[32'd162];

    assign ap_CS_fsm_state164 = ap_CS_fsm[32'd163];

    assign ap_CS_fsm_state165 = ap_CS_fsm[32'd164];

    assign ap_CS_fsm_state166 = ap_CS_fsm[32'd165];

    assign ap_CS_fsm_state167 = ap_CS_fsm[32'd166];

    assign ap_CS_fsm_state168 = ap_CS_fsm[32'd167];

    assign ap_CS_fsm_state169 = ap_CS_fsm[32'd168];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state170 = ap_CS_fsm[32'd169];

    assign ap_CS_fsm_state171 = ap_CS_fsm[32'd170];

    assign ap_CS_fsm_state172 = ap_CS_fsm[32'd171];

    assign ap_CS_fsm_state173 = ap_CS_fsm[32'd172];

    assign ap_CS_fsm_state174 = ap_CS_fsm[32'd173];

    assign ap_CS_fsm_state175 = ap_CS_fsm[32'd174];

    assign ap_CS_fsm_state176 = ap_CS_fsm[32'd175];

    assign ap_CS_fsm_state177 = ap_CS_fsm[32'd176];

    assign ap_CS_fsm_state178 = ap_CS_fsm[32'd177];

    assign ap_CS_fsm_state179 = ap_CS_fsm[32'd178];

    assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_state180 = ap_CS_fsm[32'd179];

    assign ap_CS_fsm_state181 = ap_CS_fsm[32'd180];

    assign ap_CS_fsm_state182 = ap_CS_fsm[32'd181];

    assign ap_CS_fsm_state183 = ap_CS_fsm[32'd182];

    assign ap_CS_fsm_state184 = ap_CS_fsm[32'd183];

    assign ap_CS_fsm_state185 = ap_CS_fsm[32'd184];

    assign ap_CS_fsm_state186 = ap_CS_fsm[32'd185];

    assign ap_CS_fsm_state187 = ap_CS_fsm[32'd186];

    assign ap_CS_fsm_state188 = ap_CS_fsm[32'd187];

    assign ap_CS_fsm_state189 = ap_CS_fsm[32'd188];

    assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_state190 = ap_CS_fsm[32'd189];

    assign ap_CS_fsm_state191 = ap_CS_fsm[32'd190];

    assign ap_CS_fsm_state192 = ap_CS_fsm[32'd191];

    assign ap_CS_fsm_state193 = ap_CS_fsm[32'd192];

    assign ap_CS_fsm_state194 = ap_CS_fsm[32'd193];

    assign ap_CS_fsm_state195 = ap_CS_fsm[32'd194];

    assign ap_CS_fsm_state196 = ap_CS_fsm[32'd195];

    assign ap_CS_fsm_state197 = ap_CS_fsm[32'd196];

    assign ap_CS_fsm_state198 = ap_CS_fsm[32'd197];

    assign ap_CS_fsm_state199 = ap_CS_fsm[32'd198];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_state200 = ap_CS_fsm[32'd199];

    assign ap_CS_fsm_state201 = ap_CS_fsm[32'd200];

    assign ap_CS_fsm_state202 = ap_CS_fsm[32'd201];

    assign ap_CS_fsm_state203 = ap_CS_fsm[32'd202];

    assign ap_CS_fsm_state204 = ap_CS_fsm[32'd203];

    assign ap_CS_fsm_state205 = ap_CS_fsm[32'd204];

    assign ap_CS_fsm_state206 = ap_CS_fsm[32'd205];

    assign ap_CS_fsm_state207 = ap_CS_fsm[32'd206];

    assign ap_CS_fsm_state208 = ap_CS_fsm[32'd207];

    assign ap_CS_fsm_state209 = ap_CS_fsm[32'd208];

    assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_state210 = ap_CS_fsm[32'd209];

    assign ap_CS_fsm_state211 = ap_CS_fsm[32'd210];

    assign ap_CS_fsm_state212 = ap_CS_fsm[32'd211];

    assign ap_CS_fsm_state213 = ap_CS_fsm[32'd212];

    assign ap_CS_fsm_state214 = ap_CS_fsm[32'd213];

    assign ap_CS_fsm_state215 = ap_CS_fsm[32'd214];

    assign ap_CS_fsm_state216 = ap_CS_fsm[32'd215];

    assign ap_CS_fsm_state217 = ap_CS_fsm[32'd216];

    assign ap_CS_fsm_state218 = ap_CS_fsm[32'd217];

    assign ap_CS_fsm_state219 = ap_CS_fsm[32'd218];

    assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_state220 = ap_CS_fsm[32'd219];

    assign ap_CS_fsm_state221 = ap_CS_fsm[32'd220];

    assign ap_CS_fsm_state222 = ap_CS_fsm[32'd221];

    assign ap_CS_fsm_state223 = ap_CS_fsm[32'd222];

    assign ap_CS_fsm_state224 = ap_CS_fsm[32'd223];

    assign ap_CS_fsm_state225 = ap_CS_fsm[32'd224];

    assign ap_CS_fsm_state226 = ap_CS_fsm[32'd225];

    assign ap_CS_fsm_state227 = ap_CS_fsm[32'd226];

    assign ap_CS_fsm_state228 = ap_CS_fsm[32'd227];

    assign ap_CS_fsm_state229 = ap_CS_fsm[32'd228];

    assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_state230 = ap_CS_fsm[32'd229];

    assign ap_CS_fsm_state231 = ap_CS_fsm[32'd230];

    assign ap_CS_fsm_state232 = ap_CS_fsm[32'd231];

    assign ap_CS_fsm_state233 = ap_CS_fsm[32'd232];

    assign ap_CS_fsm_state234 = ap_CS_fsm[32'd233];

    assign ap_CS_fsm_state235 = ap_CS_fsm[32'd234];

    assign ap_CS_fsm_state236 = ap_CS_fsm[32'd235];

    assign ap_CS_fsm_state237 = ap_CS_fsm[32'd236];

    assign ap_CS_fsm_state238 = ap_CS_fsm[32'd237];

    assign ap_CS_fsm_state239 = ap_CS_fsm[32'd238];

    assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_state240 = ap_CS_fsm[32'd239];

    assign ap_CS_fsm_state241 = ap_CS_fsm[32'd240];

    assign ap_CS_fsm_state242 = ap_CS_fsm[32'd241];

    assign ap_CS_fsm_state243 = ap_CS_fsm[32'd242];

    assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];

    assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];

    assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];

    assign ap_CS_fsm_state34 = ap_CS_fsm[32'd33];

    assign ap_CS_fsm_state35 = ap_CS_fsm[32'd34];

    assign ap_CS_fsm_state36 = ap_CS_fsm[32'd35];

    assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];

    assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];

    assign ap_CS_fsm_state39 = ap_CS_fsm[32'd38];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state40 = ap_CS_fsm[32'd39];

    assign ap_CS_fsm_state41 = ap_CS_fsm[32'd40];

    assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];

    assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];

    assign ap_CS_fsm_state44 = ap_CS_fsm[32'd43];

    assign ap_CS_fsm_state45 = ap_CS_fsm[32'd44];

    assign ap_CS_fsm_state46 = ap_CS_fsm[32'd45];

    assign ap_CS_fsm_state47 = ap_CS_fsm[32'd46];

    assign ap_CS_fsm_state48 = ap_CS_fsm[32'd47];

    assign ap_CS_fsm_state49 = ap_CS_fsm[32'd48];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state50 = ap_CS_fsm[32'd49];

    assign ap_CS_fsm_state51 = ap_CS_fsm[32'd50];

    assign ap_CS_fsm_state52 = ap_CS_fsm[32'd51];

    assign ap_CS_fsm_state53 = ap_CS_fsm[32'd52];

    assign ap_CS_fsm_state54 = ap_CS_fsm[32'd53];

    assign ap_CS_fsm_state55 = ap_CS_fsm[32'd54];

    assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];

    assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];

    assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];

    assign ap_CS_fsm_state59 = ap_CS_fsm[32'd58];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state60 = ap_CS_fsm[32'd59];

    assign ap_CS_fsm_state61 = ap_CS_fsm[32'd60];

    assign ap_CS_fsm_state62 = ap_CS_fsm[32'd61];

    assign ap_CS_fsm_state63 = ap_CS_fsm[32'd62];

    assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];

    assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];

    assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];

    assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];

    assign ap_CS_fsm_state68 = ap_CS_fsm[32'd67];

    assign ap_CS_fsm_state69 = ap_CS_fsm[32'd68];

    assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];

    assign ap_CS_fsm_state71 = ap_CS_fsm[32'd70];

    assign ap_CS_fsm_state72 = ap_CS_fsm[32'd71];

    assign ap_CS_fsm_state73 = ap_CS_fsm[32'd72];

    assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];

    assign ap_CS_fsm_state75 = ap_CS_fsm[32'd74];

    assign ap_CS_fsm_state76 = ap_CS_fsm[32'd75];

    assign ap_CS_fsm_state77 = ap_CS_fsm[32'd76];

    assign ap_CS_fsm_state78 = ap_CS_fsm[32'd77];

    assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

    assign ap_CS_fsm_state81 = ap_CS_fsm[32'd80];

    assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];

    assign ap_CS_fsm_state83 = ap_CS_fsm[32'd82];

    assign ap_CS_fsm_state84 = ap_CS_fsm[32'd83];

    assign ap_CS_fsm_state85 = ap_CS_fsm[32'd84];

    assign ap_CS_fsm_state86 = ap_CS_fsm[32'd85];

    assign ap_CS_fsm_state87 = ap_CS_fsm[32'd86];

    assign ap_CS_fsm_state88 = ap_CS_fsm[32'd87];

    assign ap_CS_fsm_state89 = ap_CS_fsm[32'd88];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_state90 = ap_CS_fsm[32'd89];

    assign ap_CS_fsm_state91 = ap_CS_fsm[32'd90];

    assign ap_CS_fsm_state92 = ap_CS_fsm[32'd91];

    assign ap_CS_fsm_state93 = ap_CS_fsm[32'd92];

    assign ap_CS_fsm_state94 = ap_CS_fsm[32'd93];

    assign ap_CS_fsm_state95 = ap_CS_fsm[32'd94];

    assign ap_CS_fsm_state96 = ap_CS_fsm[32'd95];

    assign ap_CS_fsm_state97 = ap_CS_fsm[32'd96];

    assign ap_CS_fsm_state98 = ap_CS_fsm[32'd97];

    assign ap_CS_fsm_state99 = ap_CS_fsm[32'd98];

    assign ap_NS_fsm_state224 = ap_NS_fsm[32'd223];

    always @(*) begin
        ap_block_state225_on_subcall_done = ((grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_done == 1'b0) | (grp_sin_or_cos_double_s_fu_421_p_done == 1'b0));
    end

    always @(*) begin
        ap_block_state79_on_subcall_done = ((grp_sin_or_cos_double_s_fu_234_ap_done == 1'b0) | (grp_sin_or_cos_double_s_fu_432_p_done == 1'b0) | (grp_sin_or_cos_double_s_fu_421_p_done == 1'b0) | (grp_atan2_cordic_double_s_fu_188_ap_done == 1'b0));
    end

    assign bitcast_ln107_fu_656_p1 = reg_427;

    assign bitcast_ln116_1_fu_761_p1 = reg_497;

    assign bitcast_ln116_fu_756_p1 = trunc_ln116_reg_1057;

    assign bitcast_ln117_1_fu_771_p1 = trunc_ln117_1_reg_1062;

    assign bitcast_ln117_fu_766_p1 = reg_501;

    assign bitcast_ln135_fu_804_p1 = reg_501;

    assign bitcast_ln137_1_fu_817_p1 = reg_530;

    assign bitcast_ln137_fu_809_p1 = trunc_ln137_reg_1122;

    assign bitcast_ln138_1_fu_831_p1 = reg_530;

    assign bitcast_ln138_fu_826_p1 = reg_497;

    assign bitcast_ln46_fu_838_p1 = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_angle_assign_3_out;

    assign bitcast_ln497_1_fu_631_p1 = t_1_fu_623_p3;

    assign bitcast_ln497_2_fu_651_p1 = t_2_fu_643_p3;

    assign bitcast_ln497_fu_610_p1 = t_fu_602_p3;

    assign data_1_fu_615_p1 = reg_419;

    assign data_2_fu_636_p1 = thetaDiff_reg_915;

    assign data_fu_594_p1 = reg_411;

    assign grp_atan2_cordic_double_s_fu_188_ap_start = grp_atan2_cordic_double_s_fu_188_ap_start_reg;

    assign grp_fu_298_p0 = $unsigned(reg_584);

    assign grp_fu_301_p0 = zext_ln57_5_fu_737_p0;

    assign grp_fu_394_p_ce = grp_fu_310_ce;

    assign grp_fu_394_p_din0 = grp_fu_310_p0;

    assign grp_fu_397_p_ce = grp_fu_319_ce;

    assign grp_fu_397_p_din0 = grp_fu_319_p0;

    assign grp_fu_397_p_din1 = grp_fu_319_p1;

    assign grp_fu_397_p_opcode = grp_fu_319_opcode;

    assign grp_fu_401_p_ce = grp_fu_323_ce;

    assign grp_fu_401_p_din0 = grp_fu_323_p0;

    assign grp_fu_401_p_din1 = grp_fu_323_p1;

    assign grp_fu_401_p_opcode = grp_fu_323_opcode;

    assign grp_fu_405_p_ce = grp_fu_333_ce;

    assign grp_fu_405_p_din0 = grp_fu_333_p0;

    assign grp_fu_405_p_din1 = grp_fu_333_p1;

    assign grp_fu_409_p_ce = 1'b1;

    assign grp_fu_409_p_din0 = grp_fu_337_p0;

    assign grp_fu_409_p_din1 = grp_fu_337_p1;

    assign grp_fu_413_p_ce = grp_fu_361_ce;

    assign grp_fu_413_p_din0 = grp_fu_361_p0;

    assign grp_fu_413_p_din1 = grp_fu_361_p1;

    assign grp_fu_413_p_opcode = grp_fu_361_opcode;

    assign grp_fu_417_p_ce = grp_fu_366_ce;

    assign grp_fu_417_p_din0 = 64'd0;

    assign grp_fu_417_p_din1 = grp_fu_366_p1;

    assign grp_fu_573_p2 = (reg_457 + 31'd12345);

    assign grp_sin_or_cos_double_s_fu_196_ap_done = grp_sin_or_cos_double_s_fu_421_p_done;

    assign grp_sin_or_cos_double_s_fu_196_ap_ready = grp_sin_or_cos_double_s_fu_421_p_ready;

    assign grp_sin_or_cos_double_s_fu_215_ap_ready = grp_sin_or_cos_double_s_fu_432_p_ready;

    assign grp_sin_or_cos_double_s_fu_234_ap_start = grp_sin_or_cos_double_s_fu_234_ap_start_reg;

    assign grp_sin_or_cos_double_s_fu_421_p_din1 = grp_sin_or_cos_double_s_fu_196_t_in;

    assign grp_sin_or_cos_double_s_fu_421_p_din2 = grp_sin_or_cos_double_s_fu_196_do_cos;

    assign grp_sin_or_cos_double_s_fu_421_p_start = grp_sin_or_cos_double_s_fu_196_ap_start_reg;

    assign grp_sin_or_cos_double_s_fu_432_p_din1 = reg_448;

    assign grp_sin_or_cos_double_s_fu_432_p_din2 = 1'd1;

    assign grp_sin_or_cos_double_s_fu_432_p_start = grp_sin_or_cos_double_s_fu_215_ap_start_reg;

    assign grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start = grp_updateMotion_Pipeline_VITIS_LOOP_45_1_fu_254_ap_start_reg;

    assign grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start = grp_updateMotion_Pipeline_VITIS_LOOP_46_2_fu_260_ap_start_reg;

    assign icmp_ln107_1_fu_680_p2 = ((trunc_ln107_fu_670_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln107_fu_674_p2 = ((tmp_fu_660_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln134_fu_778_p2 = ((i_fu_126 == 9'd500) ? 1'b1 : 1'b0);

    assign or_ln107_fu_686_p2 = (icmp_ln107_reg_926 | icmp_ln107_1_reg_931);

    assign or_ln139_7_fu_842_p4 = {
        {{bitcast_ln46_fu_838_p1}, {bitcast_ln138_1_fu_831_p1}}, {64'd0}
    };

    assign t_1_fu_623_p3 = {{1'd0}, {trunc_ln479_1_fu_619_p1}};

    assign t_2_fu_643_p3 = {{1'd0}, {trunc_ln479_2_fu_639_p1}};

    assign t_fu_602_p3 = {{1'd0}, {trunc_ln479_fu_598_p1}};

    assign tmp_fu_660_p4 = {{bitcast_ln107_fu_656_p1[62:52]}};

    assign trunc_ln107_fu_670_p1 = bitcast_ln107_fu_656_p1[51:0];

    assign trunc_ln116_fu_742_p1 = pf_q0[63:0];

    assign trunc_ln137_fu_800_p1 = pf_q0[63:0];

    assign trunc_ln479_1_fu_619_p1 = data_1_fu_615_p1[62:0];

    assign trunc_ln479_2_fu_639_p1 = data_2_fu_636_p1[62:0];

    assign trunc_ln479_fu_598_p1 = data_fu_594_p1[62:0];

    assign zext_ln134_fu_790_p1 = i_fu_126;

    assign zext_ln137_fu_821_p1 = bitcast_ln137_1_fu_817_p1;

    assign zext_ln139_fu_852_p1 = or_ln139_7_fu_842_p4;

    assign zext_ln57_1_fu_727_p1 = $unsigned(reg_579);

    assign zext_ln57_2_fu_711_p1 = $unsigned(reg_584);

    assign zext_ln57_4_fu_716_p1 = $unsigned(reg_589);

    assign zext_ln57_5_fu_737_p0 = reg_589;

    assign zext_ln57_fu_706_p1 = $unsigned(reg_579);

    always @(posedge ap_clk) begin
        pf_addr_4_reg_1117[16:9] <= 8'b00000000;
    end

endmodule  //main_updateMotion
