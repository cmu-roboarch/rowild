/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_updateSensor_Pipeline_VITIS_LOOP_173_3 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    empty_10,
    empty_11,
    empty_12,
    empty_13,
    empty,
    trunc_ln3,
    mul_ln177,
    laserReading_address0,
    laserReading_ce0,
    laserReading_q0,
    zStar_address0,
    zStar_ce0,
    zStar_q0,
    pf_load_2,
    trunc_ln188_2,
    pRand,
    bitcast_ln205,
    probability_out,
    probability_out_ap_vld,
    grp_fu_613_p_din0,
    grp_fu_613_p_dout0,
    grp_fu_613_p_ce,
    grp_fu_616_p_din0,
    grp_fu_616_p_din1,
    grp_fu_616_p_opcode,
    grp_fu_616_p_dout0,
    grp_fu_616_p_ce,
    grp_fu_597_p_din0,
    grp_fu_597_p_din1,
    grp_fu_597_p_opcode,
    grp_fu_597_p_dout0,
    grp_fu_597_p_ce,
    grp_fu_605_p_din0,
    grp_fu_605_p_din1,
    grp_fu_605_p_dout0,
    grp_fu_605_p_ce,
    grp_fu_609_p_din0,
    grp_fu_609_p_din1,
    grp_fu_609_p_dout0,
    grp_fu_609_p_ce,
    grp_fu_221_p_din0,
    grp_fu_221_p_din1,
    grp_fu_221_p_dout0,
    grp_fu_221_p_ce,
    grp_fu_620_p_din0,
    grp_fu_620_p_din1,
    grp_fu_620_p_opcode,
    grp_fu_620_p_dout0,
    grp_fu_620_p_ce,
    grp_fu_646_p_din0,
    grp_fu_646_p_din1,
    grp_fu_646_p_dout0,
    grp_fu_646_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 7'd1;
    parameter ap_ST_fsm_pp0_stage1 = 7'd2;
    parameter ap_ST_fsm_pp0_stage2 = 7'd4;
    parameter ap_ST_fsm_pp0_stage3 = 7'd8;
    parameter ap_ST_fsm_pp0_stage4 = 7'd16;
    parameter ap_ST_fsm_pp0_stage5 = 7'd32;
    parameter ap_ST_fsm_pp0_stage6 = 7'd64;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] empty_10;
    input [63:0] empty_11;
    input [63:0] empty_12;
    input [63:0] empty_13;
    input [63:0] empty;
    input [17:0] trunc_ln3;
    input [17:0] mul_ln177;
    output [17:0] laserReading_address0;
    output laserReading_ce0;
    input [31:0] laserReading_q0;
    output [7:0] zStar_address0;
    output zStar_ce0;
    input [63:0] zStar_q0;
    input [254:0] pf_load_2;
    input [51:0] trunc_ln188_2;
    input [63:0] pRand;
    input [63:0] bitcast_ln205;
    output [63:0] probability_out;
    output probability_out_ap_vld;
    output [31:0] grp_fu_613_p_din0;
    input [63:0] grp_fu_613_p_dout0;
    output grp_fu_613_p_ce;
    output [31:0] grp_fu_616_p_din0;
    output [31:0] grp_fu_616_p_din1;
    output [4:0] grp_fu_616_p_opcode;
    input [0:0] grp_fu_616_p_dout0;
    output grp_fu_616_p_ce;
    output [63:0] grp_fu_597_p_din0;
    output [63:0] grp_fu_597_p_din1;
    output [1:0] grp_fu_597_p_opcode;
    input [63:0] grp_fu_597_p_dout0;
    output grp_fu_597_p_ce;
    output [63:0] grp_fu_605_p_din0;
    output [63:0] grp_fu_605_p_din1;
    input [63:0] grp_fu_605_p_dout0;
    output grp_fu_605_p_ce;
    output [63:0] grp_fu_609_p_din0;
    output [63:0] grp_fu_609_p_din1;
    input [63:0] grp_fu_609_p_dout0;
    output grp_fu_609_p_ce;
    output [63:0] grp_fu_221_p_din0;
    output [63:0] grp_fu_221_p_din1;
    input [63:0] grp_fu_221_p_dout0;
    output grp_fu_221_p_ce;
    output [63:0] grp_fu_620_p_din0;
    output [63:0] grp_fu_620_p_din1;
    output [4:0] grp_fu_620_p_opcode;
    input [0:0] grp_fu_620_p_dout0;
    output grp_fu_620_p_ce;
    output [63:0] grp_fu_646_p_din0;
    output [63:0] grp_fu_646_p_din1;
    input [63:0] grp_fu_646_p_dout0;
    output grp_fu_646_p_ce;

    reg ap_idle;
    reg laserReading_ce0;
    reg zStar_ce0;
    reg probability_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [6:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_enable_reg_pp0_iter27;
    reg    ap_enable_reg_pp0_iter28;
    reg    ap_enable_reg_pp0_iter29;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_subdone;
    reg   [0:0] icmp_ln173_reg_655;
    reg    ap_condition_exit_pp0_iter0_stage6;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    wire   [0:0] icmp_ln173_fu_311_p2;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter1_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter2_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter3_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter4_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter5_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter6_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter7_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter8_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter9_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter10_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter11_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter12_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter13_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter14_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter15_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter16_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter17_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter18_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter19_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter20_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter21_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter22_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter23_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter24_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter25_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter26_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter27_reg;
    reg   [0:0] icmp_ln173_reg_655_pp0_iter28_reg;
    wire   [0:0] icmp_ln188_5_fu_348_p2;
    reg   [0:0] icmp_ln188_5_reg_669;
    reg   [63:0] expDist_reg_674;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    reg   [31:0] laserReading_load_reg_682;
    wire   [0:0] icmp_ln188_fu_381_p2;
    reg   [0:0] icmp_ln188_reg_689;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire   [0:0] icmp_ln188_1_fu_387_p2;
    reg   [0:0] icmp_ln188_1_reg_694;
    reg   [63:0] readDist_reg_699;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire   [0:0] and_ln188_1_fu_397_p2;
    reg   [0:0] and_ln188_1_reg_707;
    wire   [0:0] or_ln188_1_fu_441_p2;
    reg   [0:0] or_ln188_1_reg_714;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire   [0:0] and_ln188_2_fu_458_p2;
    reg   [0:0] and_ln188_2_reg_719;
    wire   [0:0] and_ln204_fu_470_p2;
    reg   [0:0] and_ln204_reg_725;
    reg   [0:0] and_ln204_reg_725_pp0_iter1_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter2_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter3_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter4_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter5_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter6_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter7_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter8_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter9_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter10_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter11_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter12_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter13_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter14_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter15_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter16_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter17_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter18_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter19_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter20_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter21_reg;
    reg   [0:0] and_ln204_reg_725_pp0_iter22_reg;
    wire   [0:0] and_ln198_fu_521_p2;
    reg   [0:0] and_ln198_reg_729;
    wire    ap_block_pp0_stage6_11001;
    reg   [0:0] and_ln198_reg_729_pp0_iter1_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter2_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter3_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter4_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter5_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter6_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter7_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter8_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter9_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter10_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter11_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter12_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter13_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter14_reg;
    reg   [0:0] and_ln198_reg_729_pp0_iter15_reg;
    wire   [63:0] trunc_ln7_fu_526_p4;
    reg   [63:0] trunc_ln7_reg_733;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter1_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter2_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter3_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter4_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter5_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter6_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter7_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter8_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter9_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter10_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter11_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter12_reg;
    reg   [63:0] trunc_ln7_reg_733_pp0_iter13_reg;
    wire   [63:0] xor_ln199_fu_535_p2;
    reg   [63:0] xor_ln199_reg_738;
    reg   [0:0] tmp_1_reg_743;
    wire   [63:0] bitcast_ln199_1_fu_541_p1;
    reg   [63:0] bitcast_ln199_1_reg_748;
    wire   [63:0] pRand_1_fu_555_p3;
    reg   [63:0] pRand_1_reg_753;
    wire   [63:0] pMax_fu_566_p3;
    reg   [63:0] pMax_reg_758;
    reg   [63:0] sub26_i_reg_763;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    reg   [63:0] sub26_i_reg_763_pp0_iter2_reg;
    reg   [63:0] mul34_i_reg_769;
    reg   [63:0] mul_i_reg_774;
    reg   [63:0] mul18_i_reg_779;
    reg   [63:0] mul41_i_reg_784;
    reg   [63:0] mul41_i_reg_784_pp0_iter3_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter4_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter5_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter6_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter7_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter8_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter9_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter10_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter11_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter12_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter13_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter14_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter15_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter16_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter17_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter18_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter19_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter20_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter21_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter22_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter23_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter24_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter25_reg;
    reg   [63:0] mul41_i_reg_784_pp0_iter26_reg;
    reg   [63:0] mul43_i_reg_789;
    reg   [63:0] mul43_i_reg_789_pp0_iter3_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter4_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter5_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter6_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter7_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter8_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter9_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter10_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter11_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter12_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter13_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter14_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter15_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter16_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter17_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter18_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter19_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter20_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter21_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter22_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter23_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter24_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter25_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter26_reg;
    reg   [63:0] mul43_i_reg_789_pp0_iter27_reg;
    reg   [63:0] mul27_i_reg_794;
    reg   [63:0] mul36_i_reg_799;
    reg   [63:0] mul36_i_reg_799_pp0_iter3_reg;
    reg   [63:0] mul36_i_reg_799_pp0_iter4_reg;
    reg   [63:0] mul36_i_reg_799_pp0_iter5_reg;
    reg   [63:0] mul36_i_reg_799_pp0_iter6_reg;
    reg   [63:0] mul31_i_reg_804;
    reg   [63:0] mul29_i_reg_809;
    wire   [63:0] grp_fu_288_p2;
    reg   [63:0] tmp_s_reg_814;
    reg   [63:0] tmp_4_reg_819;
    reg   [63:0] tmp_4_reg_819_pp0_iter6_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter7_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter8_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter9_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter10_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter11_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter12_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter13_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter14_reg;
    reg   [63:0] tmp_4_reg_819_pp0_iter15_reg;
    reg   [63:0] sub12_i_reg_824;
    reg   [63:0] div32_i_reg_829;
    reg   [63:0] n_reg_834;
    wire   [63:0] bitcast_ln199_fu_574_p1;
    reg   [63:0] pHit_reg_844;
    reg   [63:0] tmp_11_reg_849;
    reg   [63:0] mul15_i_reg_854;
    reg   [63:0] pShort_reg_859;
    reg   [63:0] mul40_i_reg_864;
    reg   [63:0] mul40_i_reg_864_pp0_iter18_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter19_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter20_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter21_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter22_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter23_reg;
    reg   [63:0] mul40_i_reg_864_pp0_iter24_reg;
    reg   [63:0] mul39_i_reg_874;
    reg   [63:0] add_i_reg_879;
    reg   [63:0] add42_i_reg_884;
    reg   [63:0] add44_i_reg_889;
    reg   [63:0] probability_1_reg_899;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage4_subdone;
    wire   [63:0] ap_phi_reg_pp0_iter0_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter1_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter2_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter3_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter4_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter5_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter6_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter7_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter8_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter9_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter10_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter11_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter12_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter13_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter14_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter15_pShort_1_reg_225;
    reg   [63:0] ap_phi_reg_pp0_iter16_pShort_1_reg_225;
    wire   [63:0] ap_phi_reg_pp0_iter0_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter1_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter2_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter3_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter4_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter5_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter6_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter7_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter8_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter9_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter10_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter11_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter12_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter13_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter14_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter15_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter16_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter17_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter18_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter19_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter20_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter21_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter22_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter23_pHit_2_reg_237;
    reg   [63:0] ap_phi_reg_pp0_iter24_pHit_2_reg_237;
    wire   [63:0] zext_ln177_fu_343_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln173_fu_326_p1;
    reg   [17:0] phi_mul_fu_114;
    wire   [17:0] add_ln174_fu_331_p2;
    wire    ap_loop_init;
    reg   [17:0] ap_sig_allocacmp_phi_mul_load;
    reg   [63:0] probability_fu_118;
    reg   [63:0] ap_sig_allocacmp_probability_load;
    wire    ap_block_pp0_stage4;
    reg   [7:0] eIdx_fu_122;
    wire   [7:0] add_ln173_fu_317_p2;
    reg   [7:0] ap_sig_allocacmp_eIdx_1;
    wire    ap_block_pp0_stage4_01001;
    wire    ap_block_pp0_stage2;
    reg   [63:0] grp_fu_257_p0;
    reg   [63:0] grp_fu_257_p1;
    wire    ap_block_pp0_stage5;
    wire    ap_block_pp0_stage1;
    wire    ap_block_pp0_stage3;
    reg   [63:0] grp_fu_262_p0;
    reg   [63:0] grp_fu_262_p1;
    wire    ap_block_pp0_stage6;
    reg   [63:0] grp_fu_267_p0;
    reg   [63:0] grp_fu_267_p1;
    reg   [63:0] grp_fu_274_p0;
    reg   [63:0] grp_fu_274_p1;
    reg   [63:0] grp_fu_279_p1;
    reg   [63:0] grp_fu_288_p1;
    wire   [17:0] add_ln177_fu_337_p2;
    wire   [31:0] bitcast_ln188_fu_364_p1;
    wire   [7:0] tmp_5_fu_367_p4;
    wire   [22:0] trunc_ln188_fu_377_p1;
    wire   [0:0] or_ln188_fu_393_p2;
    wire   [63:0] bitcast_ln188_1_fu_403_p1;
    wire   [10:0] tmp_7_fu_406_p4;
    wire   [51:0] trunc_ln188_1_fu_416_p1;
    wire   [0:0] icmp_ln188_3_fu_435_p2;
    wire   [0:0] icmp_ln188_2_fu_429_p2;
    wire   [10:0] tmp_8_fu_420_p4;
    wire   [0:0] icmp_ln188_4_fu_447_p2;
    wire   [0:0] or_ln188_2_fu_453_p2;
    wire   [0:0] and_ln204_1_fu_464_p2;
    wire   [63:0] bitcast_ln198_fu_475_p1;
    wire   [10:0] tmp_2_fu_478_p4;
    wire   [51:0] trunc_ln198_fu_488_p1;
    wire   [0:0] icmp_ln198_1_fu_498_p2;
    wire   [0:0] icmp_ln198_fu_492_p2;
    wire   [0:0] or_ln198_fu_504_p2;
    wire   [0:0] and_ln198_1_fu_510_p2;
    wire   [0:0] and_ln198_2_fu_516_p2;
    wire   [0:0] and_ln188_3_fu_545_p2;
    wire   [0:0] and_ln188_fu_550_p2;
    wire   [0:0] and_ln193_fu_562_p2;
    wire    ap_block_pp0_stage2_00001;
    reg   [1:0] grp_fu_257_opcode;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage5_00001;
    wire    ap_block_pp0_stage0_00001;
    reg   [4:0] grp_fu_279_opcode;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage6_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_condition_exit_pp0_iter28_stage4;
    reg    ap_idle_pp0_0to27;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg    ap_loop_exit_ready_pp0_iter10_reg;
    reg    ap_loop_exit_ready_pp0_iter11_reg;
    reg    ap_loop_exit_ready_pp0_iter12_reg;
    reg    ap_loop_exit_ready_pp0_iter13_reg;
    reg    ap_loop_exit_ready_pp0_iter14_reg;
    reg    ap_loop_exit_ready_pp0_iter15_reg;
    reg    ap_loop_exit_ready_pp0_iter16_reg;
    reg    ap_loop_exit_ready_pp0_iter17_reg;
    reg    ap_loop_exit_ready_pp0_iter18_reg;
    reg    ap_loop_exit_ready_pp0_iter19_reg;
    reg    ap_loop_exit_ready_pp0_iter20_reg;
    reg    ap_loop_exit_ready_pp0_iter21_reg;
    reg    ap_loop_exit_ready_pp0_iter22_reg;
    reg    ap_loop_exit_ready_pp0_iter23_reg;
    reg    ap_loop_exit_ready_pp0_iter24_reg;
    reg    ap_loop_exit_ready_pp0_iter25_reg;
    reg    ap_loop_exit_ready_pp0_iter26_reg;
    reg    ap_loop_exit_ready_pp0_iter27_reg;
    reg    ap_loop_exit_ready_pp0_iter28_reg;
    reg   [6:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to29;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    reg    ap_condition_733;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 7'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter27 = 1'b0;
        #0 ap_enable_reg_pp0_iter28 = 1'b0;
        #0 ap_enable_reg_pp0_iter29 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 phi_mul_fu_114 = 18'd0;
        #0 probability_fu_118 = 64'd0;
        #0 eIdx_fu_122 = 8'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_dexp_64ns_64ns_64_21_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(21),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dexp_64ns_64ns_64_21_full_dsp_1_U178 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd0),
        .din1(grp_fu_288_p1),
        .ce(1'b1),
        .dout(grp_fu_288_p2)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage6),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (ap_loop_exit_ready_pp0_iter28_reg == 1'b1) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage6)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter27 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter28 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter29 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter29 == 1'b1))) begin
                ap_enable_reg_pp0_iter29 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter17_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter17_reg <= ap_loop_exit_ready_pp0_iter16_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter18_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter18_reg <= ap_loop_exit_ready_pp0_iter17_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter19_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter19_reg <= ap_loop_exit_ready_pp0_iter18_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter20_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter20_reg <= ap_loop_exit_ready_pp0_iter19_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter21_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter21_reg <= ap_loop_exit_ready_pp0_iter20_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter22_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter22_reg <= ap_loop_exit_ready_pp0_iter21_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter23_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter23_reg <= ap_loop_exit_ready_pp0_iter22_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter24_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter24_reg <= ap_loop_exit_ready_pp0_iter23_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter25_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter25_reg <= ap_loop_exit_ready_pp0_iter24_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter26_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter26_reg <= ap_loop_exit_ready_pp0_iter25_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter27_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter27_reg <= ap_loop_exit_ready_pp0_iter26_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter28_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter28_reg <= ap_loop_exit_ready_pp0_iter27_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter16 == 1'b1) & (icmp_ln173_reg_655_pp0_iter16_reg == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'd1 == and_ln198_reg_729_pp0_iter15_reg) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            ap_phi_reg_pp0_iter16_pShort_1_reg_225 <= pShort_reg_859;
        end else if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter16_pShort_1_reg_225 <= ap_phi_reg_pp0_iter15_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_condition_733)) begin
            if (((1'd0 == and_ln204_reg_725) & (icmp_ln173_reg_655 == 1'd0))) begin
                ap_phi_reg_pp0_iter1_pHit_2_reg_237 <= 64'd0;
            end else if ((1'b1 == 1'b1)) begin
                ap_phi_reg_pp0_iter1_pHit_2_reg_237 <= ap_phi_reg_pp0_iter0_pHit_2_reg_237;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'd0 == and_ln198_reg_729) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_pShort_1_reg_225 <= 64'd0;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter1_pShort_1_reg_225 <= ap_phi_reg_pp0_iter0_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter23 == 1'b1) & (icmp_ln173_reg_655_pp0_iter23_reg == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'd1 == and_ln204_reg_725_pp0_iter22_reg) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            ap_phi_reg_pp0_iter23_pHit_2_reg_237 <= grp_fu_221_p_dout0;
        end else if (((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter23_pHit_2_reg_237 <= ap_phi_reg_pp0_iter22_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            if (((icmp_ln173_fu_311_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                eIdx_fu_122 <= add_ln173_fu_317_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                eIdx_fu_122 <= 8'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            if (((icmp_ln173_fu_311_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                phi_mul_fu_114 <= add_ln174_fu_331_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                phi_mul_fu_114 <= 18'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            probability_fu_118 <= 64'd4607182418800017408;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter29 == 1'b1))) begin
            probability_fu_118 <= probability_1_reg_899;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter27 == 1'b1))) begin
            add42_i_reg_884 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter28 == 1'b1))) begin
            add44_i_reg_889 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            add_i_reg_879 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            and_ln188_1_reg_707 <= and_ln188_1_fu_397_p2;
            mul40_i_reg_864_pp0_iter18_reg <= mul40_i_reg_864;
            mul40_i_reg_864_pp0_iter19_reg <= mul40_i_reg_864_pp0_iter18_reg;
            mul40_i_reg_864_pp0_iter20_reg <= mul40_i_reg_864_pp0_iter19_reg;
            mul40_i_reg_864_pp0_iter21_reg <= mul40_i_reg_864_pp0_iter20_reg;
            mul40_i_reg_864_pp0_iter22_reg <= mul40_i_reg_864_pp0_iter21_reg;
            mul40_i_reg_864_pp0_iter23_reg <= mul40_i_reg_864_pp0_iter22_reg;
            mul40_i_reg_864_pp0_iter24_reg <= mul40_i_reg_864_pp0_iter23_reg;
            readDist_reg_699 <= grp_fu_613_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5_11001))) begin
            and_ln188_2_reg_719 <= and_ln188_2_fu_458_p2;
            and_ln204_reg_725 <= and_ln204_fu_470_p2;
            and_ln204_reg_725_pp0_iter10_reg <= and_ln204_reg_725_pp0_iter9_reg;
            and_ln204_reg_725_pp0_iter11_reg <= and_ln204_reg_725_pp0_iter10_reg;
            and_ln204_reg_725_pp0_iter12_reg <= and_ln204_reg_725_pp0_iter11_reg;
            and_ln204_reg_725_pp0_iter13_reg <= and_ln204_reg_725_pp0_iter12_reg;
            and_ln204_reg_725_pp0_iter14_reg <= and_ln204_reg_725_pp0_iter13_reg;
            and_ln204_reg_725_pp0_iter15_reg <= and_ln204_reg_725_pp0_iter14_reg;
            and_ln204_reg_725_pp0_iter16_reg <= and_ln204_reg_725_pp0_iter15_reg;
            and_ln204_reg_725_pp0_iter17_reg <= and_ln204_reg_725_pp0_iter16_reg;
            and_ln204_reg_725_pp0_iter18_reg <= and_ln204_reg_725_pp0_iter17_reg;
            and_ln204_reg_725_pp0_iter19_reg <= and_ln204_reg_725_pp0_iter18_reg;
            and_ln204_reg_725_pp0_iter1_reg <= and_ln204_reg_725;
            and_ln204_reg_725_pp0_iter20_reg <= and_ln204_reg_725_pp0_iter19_reg;
            and_ln204_reg_725_pp0_iter21_reg <= and_ln204_reg_725_pp0_iter20_reg;
            and_ln204_reg_725_pp0_iter22_reg <= and_ln204_reg_725_pp0_iter21_reg;
            and_ln204_reg_725_pp0_iter2_reg <= and_ln204_reg_725_pp0_iter1_reg;
            and_ln204_reg_725_pp0_iter3_reg <= and_ln204_reg_725_pp0_iter2_reg;
            and_ln204_reg_725_pp0_iter4_reg <= and_ln204_reg_725_pp0_iter3_reg;
            and_ln204_reg_725_pp0_iter5_reg <= and_ln204_reg_725_pp0_iter4_reg;
            and_ln204_reg_725_pp0_iter6_reg <= and_ln204_reg_725_pp0_iter5_reg;
            and_ln204_reg_725_pp0_iter7_reg <= and_ln204_reg_725_pp0_iter6_reg;
            and_ln204_reg_725_pp0_iter8_reg <= and_ln204_reg_725_pp0_iter7_reg;
            and_ln204_reg_725_pp0_iter9_reg <= and_ln204_reg_725_pp0_iter8_reg;
            or_ln188_1_reg_714 <= or_ln188_1_fu_441_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            and_ln198_reg_729 <= and_ln198_fu_521_p2;
            and_ln198_reg_729_pp0_iter10_reg <= and_ln198_reg_729_pp0_iter9_reg;
            and_ln198_reg_729_pp0_iter11_reg <= and_ln198_reg_729_pp0_iter10_reg;
            and_ln198_reg_729_pp0_iter12_reg <= and_ln198_reg_729_pp0_iter11_reg;
            and_ln198_reg_729_pp0_iter13_reg <= and_ln198_reg_729_pp0_iter12_reg;
            and_ln198_reg_729_pp0_iter14_reg <= and_ln198_reg_729_pp0_iter13_reg;
            and_ln198_reg_729_pp0_iter15_reg <= and_ln198_reg_729_pp0_iter14_reg;
            and_ln198_reg_729_pp0_iter1_reg <= and_ln198_reg_729;
            and_ln198_reg_729_pp0_iter2_reg <= and_ln198_reg_729_pp0_iter1_reg;
            and_ln198_reg_729_pp0_iter3_reg <= and_ln198_reg_729_pp0_iter2_reg;
            and_ln198_reg_729_pp0_iter4_reg <= and_ln198_reg_729_pp0_iter3_reg;
            and_ln198_reg_729_pp0_iter5_reg <= and_ln198_reg_729_pp0_iter4_reg;
            and_ln198_reg_729_pp0_iter6_reg <= and_ln198_reg_729_pp0_iter5_reg;
            and_ln198_reg_729_pp0_iter7_reg <= and_ln198_reg_729_pp0_iter6_reg;
            and_ln198_reg_729_pp0_iter8_reg <= and_ln198_reg_729_pp0_iter7_reg;
            and_ln198_reg_729_pp0_iter9_reg <= and_ln198_reg_729_pp0_iter8_reg;
            mul36_i_reg_799_pp0_iter3_reg <= mul36_i_reg_799;
            mul36_i_reg_799_pp0_iter4_reg <= mul36_i_reg_799_pp0_iter3_reg;
            mul36_i_reg_799_pp0_iter5_reg <= mul36_i_reg_799_pp0_iter4_reg;
            mul36_i_reg_799_pp0_iter6_reg <= mul36_i_reg_799_pp0_iter5_reg;
            trunc_ln7_reg_733 <= {{pf_load_2[127:64]}};
            trunc_ln7_reg_733_pp0_iter10_reg <= trunc_ln7_reg_733_pp0_iter9_reg;
            trunc_ln7_reg_733_pp0_iter11_reg <= trunc_ln7_reg_733_pp0_iter10_reg;
            trunc_ln7_reg_733_pp0_iter12_reg <= trunc_ln7_reg_733_pp0_iter11_reg;
            trunc_ln7_reg_733_pp0_iter13_reg <= trunc_ln7_reg_733_pp0_iter12_reg;
            trunc_ln7_reg_733_pp0_iter1_reg <= trunc_ln7_reg_733;
            trunc_ln7_reg_733_pp0_iter2_reg <= trunc_ln7_reg_733_pp0_iter1_reg;
            trunc_ln7_reg_733_pp0_iter3_reg <= trunc_ln7_reg_733_pp0_iter2_reg;
            trunc_ln7_reg_733_pp0_iter4_reg <= trunc_ln7_reg_733_pp0_iter3_reg;
            trunc_ln7_reg_733_pp0_iter5_reg <= trunc_ln7_reg_733_pp0_iter4_reg;
            trunc_ln7_reg_733_pp0_iter6_reg <= trunc_ln7_reg_733_pp0_iter5_reg;
            trunc_ln7_reg_733_pp0_iter7_reg <= trunc_ln7_reg_733_pp0_iter6_reg;
            trunc_ln7_reg_733_pp0_iter8_reg <= trunc_ln7_reg_733_pp0_iter7_reg;
            trunc_ln7_reg_733_pp0_iter9_reg <= trunc_ln7_reg_733_pp0_iter8_reg;
            xor_ln199_reg_738 <= xor_ln199_fu_535_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter10_pHit_2_reg_237   <= ap_phi_reg_pp0_iter9_pHit_2_reg_237;
            ap_phi_reg_pp0_iter10_pShort_1_reg_225 <= ap_phi_reg_pp0_iter9_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter11_pHit_2_reg_237   <= ap_phi_reg_pp0_iter10_pHit_2_reg_237;
            ap_phi_reg_pp0_iter11_pShort_1_reg_225 <= ap_phi_reg_pp0_iter10_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter12_pHit_2_reg_237   <= ap_phi_reg_pp0_iter11_pHit_2_reg_237;
            ap_phi_reg_pp0_iter12_pShort_1_reg_225 <= ap_phi_reg_pp0_iter11_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter13_pHit_2_reg_237   <= ap_phi_reg_pp0_iter12_pHit_2_reg_237;
            ap_phi_reg_pp0_iter13_pShort_1_reg_225 <= ap_phi_reg_pp0_iter12_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter14_pHit_2_reg_237   <= ap_phi_reg_pp0_iter13_pHit_2_reg_237;
            ap_phi_reg_pp0_iter14_pShort_1_reg_225 <= ap_phi_reg_pp0_iter13_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter15_pHit_2_reg_237   <= ap_phi_reg_pp0_iter14_pHit_2_reg_237;
            ap_phi_reg_pp0_iter15_pShort_1_reg_225 <= ap_phi_reg_pp0_iter14_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter16_pHit_2_reg_237 <= ap_phi_reg_pp0_iter15_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter17_pHit_2_reg_237 <= ap_phi_reg_pp0_iter16_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter18_pHit_2_reg_237 <= ap_phi_reg_pp0_iter17_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter18 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter19_pHit_2_reg_237 <= ap_phi_reg_pp0_iter18_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter20_pHit_2_reg_237 <= ap_phi_reg_pp0_iter19_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter20 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter21_pHit_2_reg_237 <= ap_phi_reg_pp0_iter20_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter22_pHit_2_reg_237 <= ap_phi_reg_pp0_iter21_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter23 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter24_pHit_2_reg_237 <= ap_phi_reg_pp0_iter23_pHit_2_reg_237;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter2_pHit_2_reg_237 <= ap_phi_reg_pp0_iter1_pHit_2_reg_237;
            ap_phi_reg_pp0_iter2_pShort_1_reg_225 <= ap_phi_reg_pp0_iter1_pShort_1_reg_225;
            mul_i_reg_774 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter3_pHit_2_reg_237 <= ap_phi_reg_pp0_iter2_pHit_2_reg_237;
            ap_phi_reg_pp0_iter3_pShort_1_reg_225 <= ap_phi_reg_pp0_iter2_pShort_1_reg_225;
            mul36_i_reg_799 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter4_pHit_2_reg_237   <= ap_phi_reg_pp0_iter3_pHit_2_reg_237;
            ap_phi_reg_pp0_iter4_pShort_1_reg_225 <= ap_phi_reg_pp0_iter3_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter5_pHit_2_reg_237 <= ap_phi_reg_pp0_iter4_pHit_2_reg_237;
            ap_phi_reg_pp0_iter5_pShort_1_reg_225 <= ap_phi_reg_pp0_iter4_pShort_1_reg_225;
            tmp_s_reg_814 <= grp_fu_288_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter6_pHit_2_reg_237 <= ap_phi_reg_pp0_iter5_pHit_2_reg_237;
            ap_phi_reg_pp0_iter6_pShort_1_reg_225 <= ap_phi_reg_pp0_iter5_pShort_1_reg_225;
            sub12_i_reg_824 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter7_pHit_2_reg_237   <= ap_phi_reg_pp0_iter6_pHit_2_reg_237;
            ap_phi_reg_pp0_iter7_pShort_1_reg_225 <= ap_phi_reg_pp0_iter6_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter8_pHit_2_reg_237   <= ap_phi_reg_pp0_iter7_pHit_2_reg_237;
            ap_phi_reg_pp0_iter8_pShort_1_reg_225 <= ap_phi_reg_pp0_iter7_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001))) begin
            ap_phi_reg_pp0_iter9_pHit_2_reg_237   <= ap_phi_reg_pp0_iter8_pHit_2_reg_237;
            ap_phi_reg_pp0_iter9_pShort_1_reg_225 <= ap_phi_reg_pp0_iter8_pShort_1_reg_225;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            bitcast_ln199_1_reg_748 <= bitcast_ln199_1_fu_541_p1;
            icmp_ln173_reg_655 <= icmp_ln173_fu_311_p2;
            icmp_ln173_reg_655_pp0_iter10_reg <= icmp_ln173_reg_655_pp0_iter9_reg;
            icmp_ln173_reg_655_pp0_iter11_reg <= icmp_ln173_reg_655_pp0_iter10_reg;
            icmp_ln173_reg_655_pp0_iter12_reg <= icmp_ln173_reg_655_pp0_iter11_reg;
            icmp_ln173_reg_655_pp0_iter13_reg <= icmp_ln173_reg_655_pp0_iter12_reg;
            icmp_ln173_reg_655_pp0_iter14_reg <= icmp_ln173_reg_655_pp0_iter13_reg;
            icmp_ln173_reg_655_pp0_iter15_reg <= icmp_ln173_reg_655_pp0_iter14_reg;
            icmp_ln173_reg_655_pp0_iter16_reg <= icmp_ln173_reg_655_pp0_iter15_reg;
            icmp_ln173_reg_655_pp0_iter17_reg <= icmp_ln173_reg_655_pp0_iter16_reg;
            icmp_ln173_reg_655_pp0_iter18_reg <= icmp_ln173_reg_655_pp0_iter17_reg;
            icmp_ln173_reg_655_pp0_iter19_reg <= icmp_ln173_reg_655_pp0_iter18_reg;
            icmp_ln173_reg_655_pp0_iter1_reg <= icmp_ln173_reg_655;
            icmp_ln173_reg_655_pp0_iter20_reg <= icmp_ln173_reg_655_pp0_iter19_reg;
            icmp_ln173_reg_655_pp0_iter21_reg <= icmp_ln173_reg_655_pp0_iter20_reg;
            icmp_ln173_reg_655_pp0_iter22_reg <= icmp_ln173_reg_655_pp0_iter21_reg;
            icmp_ln173_reg_655_pp0_iter23_reg <= icmp_ln173_reg_655_pp0_iter22_reg;
            icmp_ln173_reg_655_pp0_iter24_reg <= icmp_ln173_reg_655_pp0_iter23_reg;
            icmp_ln173_reg_655_pp0_iter25_reg <= icmp_ln173_reg_655_pp0_iter24_reg;
            icmp_ln173_reg_655_pp0_iter26_reg <= icmp_ln173_reg_655_pp0_iter25_reg;
            icmp_ln173_reg_655_pp0_iter27_reg <= icmp_ln173_reg_655_pp0_iter26_reg;
            icmp_ln173_reg_655_pp0_iter28_reg <= icmp_ln173_reg_655_pp0_iter27_reg;
            icmp_ln173_reg_655_pp0_iter2_reg <= icmp_ln173_reg_655_pp0_iter1_reg;
            icmp_ln173_reg_655_pp0_iter3_reg <= icmp_ln173_reg_655_pp0_iter2_reg;
            icmp_ln173_reg_655_pp0_iter4_reg <= icmp_ln173_reg_655_pp0_iter3_reg;
            icmp_ln173_reg_655_pp0_iter5_reg <= icmp_ln173_reg_655_pp0_iter4_reg;
            icmp_ln173_reg_655_pp0_iter6_reg <= icmp_ln173_reg_655_pp0_iter5_reg;
            icmp_ln173_reg_655_pp0_iter7_reg <= icmp_ln173_reg_655_pp0_iter6_reg;
            icmp_ln173_reg_655_pp0_iter8_reg <= icmp_ln173_reg_655_pp0_iter7_reg;
            icmp_ln173_reg_655_pp0_iter9_reg <= icmp_ln173_reg_655_pp0_iter8_reg;
            icmp_ln188_5_reg_669 <= icmp_ln188_5_fu_348_p2;
            tmp_4_reg_819_pp0_iter10_reg <= tmp_4_reg_819_pp0_iter9_reg;
            tmp_4_reg_819_pp0_iter11_reg <= tmp_4_reg_819_pp0_iter10_reg;
            tmp_4_reg_819_pp0_iter12_reg <= tmp_4_reg_819_pp0_iter11_reg;
            tmp_4_reg_819_pp0_iter13_reg <= tmp_4_reg_819_pp0_iter12_reg;
            tmp_4_reg_819_pp0_iter14_reg <= tmp_4_reg_819_pp0_iter13_reg;
            tmp_4_reg_819_pp0_iter15_reg <= tmp_4_reg_819_pp0_iter14_reg;
            tmp_4_reg_819_pp0_iter6_reg <= tmp_4_reg_819;
            tmp_4_reg_819_pp0_iter7_reg <= tmp_4_reg_819_pp0_iter6_reg;
            tmp_4_reg_819_pp0_iter8_reg <= tmp_4_reg_819_pp0_iter7_reg;
            tmp_4_reg_819_pp0_iter9_reg <= tmp_4_reg_819_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            div32_i_reg_829 <= grp_fu_221_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            expDist_reg_674 <= zStar_q0;
            laserReading_load_reg_682 <= laserReading_q0;
            mul41_i_reg_784_pp0_iter10_reg <= mul41_i_reg_784_pp0_iter9_reg;
            mul41_i_reg_784_pp0_iter11_reg <= mul41_i_reg_784_pp0_iter10_reg;
            mul41_i_reg_784_pp0_iter12_reg <= mul41_i_reg_784_pp0_iter11_reg;
            mul41_i_reg_784_pp0_iter13_reg <= mul41_i_reg_784_pp0_iter12_reg;
            mul41_i_reg_784_pp0_iter14_reg <= mul41_i_reg_784_pp0_iter13_reg;
            mul41_i_reg_784_pp0_iter15_reg <= mul41_i_reg_784_pp0_iter14_reg;
            mul41_i_reg_784_pp0_iter16_reg <= mul41_i_reg_784_pp0_iter15_reg;
            mul41_i_reg_784_pp0_iter17_reg <= mul41_i_reg_784_pp0_iter16_reg;
            mul41_i_reg_784_pp0_iter18_reg <= mul41_i_reg_784_pp0_iter17_reg;
            mul41_i_reg_784_pp0_iter19_reg <= mul41_i_reg_784_pp0_iter18_reg;
            mul41_i_reg_784_pp0_iter20_reg <= mul41_i_reg_784_pp0_iter19_reg;
            mul41_i_reg_784_pp0_iter21_reg <= mul41_i_reg_784_pp0_iter20_reg;
            mul41_i_reg_784_pp0_iter22_reg <= mul41_i_reg_784_pp0_iter21_reg;
            mul41_i_reg_784_pp0_iter23_reg <= mul41_i_reg_784_pp0_iter22_reg;
            mul41_i_reg_784_pp0_iter24_reg <= mul41_i_reg_784_pp0_iter23_reg;
            mul41_i_reg_784_pp0_iter25_reg <= mul41_i_reg_784_pp0_iter24_reg;
            mul41_i_reg_784_pp0_iter26_reg <= mul41_i_reg_784_pp0_iter25_reg;
            mul41_i_reg_784_pp0_iter3_reg <= mul41_i_reg_784;
            mul41_i_reg_784_pp0_iter4_reg <= mul41_i_reg_784_pp0_iter3_reg;
            mul41_i_reg_784_pp0_iter5_reg <= mul41_i_reg_784_pp0_iter4_reg;
            mul41_i_reg_784_pp0_iter6_reg <= mul41_i_reg_784_pp0_iter5_reg;
            mul41_i_reg_784_pp0_iter7_reg <= mul41_i_reg_784_pp0_iter6_reg;
            mul41_i_reg_784_pp0_iter8_reg <= mul41_i_reg_784_pp0_iter7_reg;
            mul41_i_reg_784_pp0_iter9_reg <= mul41_i_reg_784_pp0_iter8_reg;
            mul43_i_reg_789_pp0_iter10_reg <= mul43_i_reg_789_pp0_iter9_reg;
            mul43_i_reg_789_pp0_iter11_reg <= mul43_i_reg_789_pp0_iter10_reg;
            mul43_i_reg_789_pp0_iter12_reg <= mul43_i_reg_789_pp0_iter11_reg;
            mul43_i_reg_789_pp0_iter13_reg <= mul43_i_reg_789_pp0_iter12_reg;
            mul43_i_reg_789_pp0_iter14_reg <= mul43_i_reg_789_pp0_iter13_reg;
            mul43_i_reg_789_pp0_iter15_reg <= mul43_i_reg_789_pp0_iter14_reg;
            mul43_i_reg_789_pp0_iter16_reg <= mul43_i_reg_789_pp0_iter15_reg;
            mul43_i_reg_789_pp0_iter17_reg <= mul43_i_reg_789_pp0_iter16_reg;
            mul43_i_reg_789_pp0_iter18_reg <= mul43_i_reg_789_pp0_iter17_reg;
            mul43_i_reg_789_pp0_iter19_reg <= mul43_i_reg_789_pp0_iter18_reg;
            mul43_i_reg_789_pp0_iter20_reg <= mul43_i_reg_789_pp0_iter19_reg;
            mul43_i_reg_789_pp0_iter21_reg <= mul43_i_reg_789_pp0_iter20_reg;
            mul43_i_reg_789_pp0_iter22_reg <= mul43_i_reg_789_pp0_iter21_reg;
            mul43_i_reg_789_pp0_iter23_reg <= mul43_i_reg_789_pp0_iter22_reg;
            mul43_i_reg_789_pp0_iter24_reg <= mul43_i_reg_789_pp0_iter23_reg;
            mul43_i_reg_789_pp0_iter25_reg <= mul43_i_reg_789_pp0_iter24_reg;
            mul43_i_reg_789_pp0_iter26_reg <= mul43_i_reg_789_pp0_iter25_reg;
            mul43_i_reg_789_pp0_iter27_reg <= mul43_i_reg_789_pp0_iter26_reg;
            mul43_i_reg_789_pp0_iter3_reg <= mul43_i_reg_789;
            mul43_i_reg_789_pp0_iter4_reg <= mul43_i_reg_789_pp0_iter3_reg;
            mul43_i_reg_789_pp0_iter5_reg <= mul43_i_reg_789_pp0_iter4_reg;
            mul43_i_reg_789_pp0_iter6_reg <= mul43_i_reg_789_pp0_iter5_reg;
            mul43_i_reg_789_pp0_iter7_reg <= mul43_i_reg_789_pp0_iter6_reg;
            mul43_i_reg_789_pp0_iter8_reg <= mul43_i_reg_789_pp0_iter7_reg;
            mul43_i_reg_789_pp0_iter9_reg <= mul43_i_reg_789_pp0_iter8_reg;
            pMax_reg_758[61 : 52] <= pMax_fu_566_p3[61 : 52];
            pRand_1_reg_753 <= pRand_1_fu_555_p3;
            tmp_11_reg_849 <= grp_fu_646_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            icmp_ln188_1_reg_694 <= icmp_ln188_1_fu_387_p2;
            icmp_ln188_reg_689   <= icmp_ln188_fu_381_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            mul15_i_reg_854 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            mul18_i_reg_779 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            mul27_i_reg_794 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5_11001))) begin
            mul29_i_reg_809 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            mul31_i_reg_804 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5_11001))) begin
            mul34_i_reg_769 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter25 == 1'b1))) begin
            mul39_i_reg_874 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001))) begin
            mul40_i_reg_864 <= grp_fu_605_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            mul41_i_reg_784 <= grp_fu_605_p_dout0;
            mul43_i_reg_789 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            n_reg_834 <= grp_fu_221_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            pHit_reg_844 <= grp_fu_288_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_11001))) begin
            pShort_reg_859 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter29 == 1'b1))) begin
            probability_1_reg_899 <= grp_fu_609_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            sub26_i_reg_763 <= grp_fu_597_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            sub26_i_reg_763_pp0_iter2_reg <= sub26_i_reg_763;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            tmp_1_reg_743 <= grp_fu_620_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            tmp_4_reg_819 <= grp_fu_288_p2;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (icmp_ln173_reg_655 == 1'd1) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
            ap_condition_exit_pp0_iter0_stage6 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage6 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln173_reg_655_pp0_iter28_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter28 == 1'b1))) begin
            ap_condition_exit_pp0_iter28_stage4 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter28_stage4 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage4) & (ap_loop_exit_ready_pp0_iter28_reg == 1'b1) & (1'b0 == ap_block_pp0_stage4_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0) 
    & (ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0) & (ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0))) begin
            ap_idle_pp0_0to27 = 1'b1;
        end else begin
            ap_idle_pp0_0to27 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0) & (ap_enable_reg_pp0_iter26 == 1'b0) 
    & (ap_enable_reg_pp0_iter25 == 1'b0))) begin
            ap_idle_pp0_1to29 = 1'b1;
        end else begin
            ap_idle_pp0_1to29 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_eIdx_1 = 8'd0;
        end else begin
            ap_sig_allocacmp_eIdx_1 = eIdx_fu_122;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_phi_mul_load = 18'd0;
        end else begin
            ap_sig_allocacmp_phi_mul_load = phi_mul_fu_114;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter29 == 1'b1))) begin
            ap_sig_allocacmp_probability_load = probability_1_reg_899;
        end else begin
            ap_sig_allocacmp_probability_load = probability_fu_118;
        end
    end

    always @(*) begin
        if ((((ap_enable_reg_pp0_iter5 == 1'b1) & (icmp_ln173_reg_655_pp0_iter4_reg == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'd1 == and_ln198_reg_729_pp0_iter4_reg) & (1'b0 == ap_block_pp0_stage0_00001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'd1 == and_ln204_fu_470_p2) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage5_00001)))) begin
            grp_fu_257_opcode = 2'd1;
        end else if ((((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter27 == 1'b1)) | ((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter26 == 1'b1)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter25 == 1'b1)))) begin
            grp_fu_257_opcode = 2'd0;
        end else begin
            grp_fu_257_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter27 == 1'b1))) begin
            grp_fu_257_p0 = add42_i_reg_884;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            grp_fu_257_p0 = add_i_reg_879;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter25 == 1'b1))) begin
            grp_fu_257_p0 = mul39_i_reg_874;
        end else if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_257_p0 = 64'd4607182418800017408;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_257_p0 = readDist_reg_699;
        end else begin
            grp_fu_257_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter27 == 1'b1))) begin
            grp_fu_257_p1 = mul43_i_reg_789_pp0_iter27_reg;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter26 == 1'b1))) begin
            grp_fu_257_p1 = mul41_i_reg_784_pp0_iter26_reg;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter25 == 1'b1))) begin
            grp_fu_257_p1 = mul40_i_reg_864_pp0_iter24_reg;
        end else if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_257_p1 = tmp_s_reg_814;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_257_p1 = expDist_reg_674;
        end else begin
            grp_fu_257_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_262_p0 = empty_11;
        end else if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_262_p0 = n_reg_834;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_262_p0 = sub26_i_reg_763;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_262_p0 = empty_12;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_262_p0 = readDist_reg_699;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_262_p0 = expDist_reg_674;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_262_p0 = bitcast_ln205;
        end else begin
            grp_fu_262_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4))) begin
            grp_fu_262_p1 = ap_phi_reg_pp0_iter16_pShort_1_reg_225;
        end else if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_262_p1 = bitcast_ln199_fu_574_p1;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_262_p1 = 64'd13826050856027422720;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_262_p1 = pMax_reg_758;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_262_p1 = bitcast_ln199_1_reg_748;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_262_p1 = bitcast_ln199_1_fu_541_p1;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_262_p1 = 64'd4618760256180340048;
        end else begin
            grp_fu_262_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter28 == 1'b1))) begin
            grp_fu_267_p0 = ap_sig_allocacmp_probability_load;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_267_p0 = empty_10;
        end else if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_267_p0 = mul15_i_reg_854;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_267_p0 = mul27_i_reg_794;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_267_p0 = bitcast_ln205;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_267_p0 = mul34_i_reg_769;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_267_p0 = empty_13;
        end else begin
            grp_fu_267_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter28 == 1'b1))) begin
            grp_fu_267_p1 = add44_i_reg_889;
        end else if (((ap_enable_reg_pp0_iter24 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_267_p1 = ap_phi_reg_pp0_iter24_pHit_2_reg_237;
        end else if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (1'b0 == ap_block_pp0_stage3))) begin
            grp_fu_267_p1 = tmp_4_reg_819_pp0_iter15_reg;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_267_p1 = sub26_i_reg_763_pp0_iter2_reg;
        end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)))) begin
            grp_fu_267_p1 = bitcast_ln205;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_267_p1 = pRand_1_reg_753;
        end else begin
            grp_fu_267_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_274_p0 = pHit_reg_844;
        end else if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_274_p0 = 64'd4607182418800017408;
        end else if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_274_p0 = mul29_i_reg_809;
        end else begin
            grp_fu_274_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_274_p1 = tmp_11_reg_849;
        end else if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_274_p1 = sub12_i_reg_824;
        end else if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6))) begin
            grp_fu_274_p1 = mul31_i_reg_804;
        end else begin
            grp_fu_274_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage0_00001))) begin
            grp_fu_279_opcode = 5'd4;
        end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage6_00001))) begin
            grp_fu_279_opcode = 5'd3;
        end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage4_00001)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (icmp_ln173_reg_655 == 1'd0) & (1'b0 == ap_block_pp0_stage5_00001)))) begin
            grp_fu_279_opcode = 5'd5;
        end else begin
            grp_fu_279_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5) & (1'b0 == ap_block_pp0_stage5))) begin
            grp_fu_279_p1 = expDist_reg_674;
        end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6)))) begin
            grp_fu_279_p1 = empty;
        end else begin
            grp_fu_279_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (1'b0 == ap_block_pp0_stage2))) begin
            grp_fu_288_p1 = div32_i_reg_829;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            grp_fu_288_p1 = mul18_i_reg_779;
        end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            grp_fu_288_p1 = mul_i_reg_774;
        end else begin
            grp_fu_288_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            laserReading_ce0 = 1'b1;
        end else begin
            laserReading_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln173_reg_655_pp0_iter28_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (1'b0 == ap_block_pp0_stage4_11001))) begin
            probability_out_ap_vld = 1'b1;
        end else begin
            probability_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            zStar_ce0 = 1'b1;
        end else begin
            zStar_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to29 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if (((1'b1 == ap_condition_exit_pp0_iter28_stage4) & (ap_idle_pp0_0to27 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln173_fu_317_p2 = (ap_sig_allocacmp_eIdx_1 + 8'd1);

    assign add_ln174_fu_331_p2 = (ap_sig_allocacmp_phi_mul_load + trunc_ln3);

    assign add_ln177_fu_337_p2 = (mul_ln177 + ap_sig_allocacmp_phi_mul_load);

    assign and_ln188_1_fu_397_p2 = (or_ln188_fu_393_p2 & grp_fu_616_p_dout0);

    assign and_ln188_2_fu_458_p2 = (or_ln188_2_fu_453_p2 & or_ln188_1_fu_441_p2);

    assign and_ln188_3_fu_545_p2 = (grp_fu_620_p_dout0 & and_ln188_2_reg_719);

    assign and_ln188_fu_550_p2 = (and_ln188_3_fu_545_p2 & and_ln188_1_reg_707);

    assign and_ln193_fu_562_p2 = (tmp_1_reg_743 & and_ln188_2_reg_719);

    assign and_ln198_1_fu_510_p2 = (or_ln198_fu_504_p2 & grp_fu_620_p_dout0);

    assign and_ln198_2_fu_516_p2 = (or_ln188_1_reg_714 & and_ln198_1_fu_510_p2);

    assign and_ln198_fu_521_p2 = (and_ln198_2_fu_516_p2 & and_ln188_1_reg_707);

    assign and_ln204_1_fu_464_p2 = (grp_fu_620_p_dout0 & and_ln188_2_fu_458_p2);

    assign and_ln204_fu_470_p2 = (and_ln204_1_fu_464_p2 & and_ln188_1_reg_707);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    always @(*) begin
        ap_condition_733 = ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6) & (1'b0 == ap_block_pp0_stage6_11001));
    end

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage6;

    assign ap_phi_reg_pp0_iter0_pHit_2_reg_237 = 'bx;

    assign ap_phi_reg_pp0_iter0_pShort_1_reg_225 = 'bx;

    assign bitcast_ln188_1_fu_403_p1 = readDist_reg_699;

    assign bitcast_ln188_fu_364_p1 = laserReading_load_reg_682;

    assign bitcast_ln198_fu_475_p1 = expDist_reg_674;

    assign bitcast_ln199_1_fu_541_p1 = xor_ln199_reg_738;

    assign bitcast_ln199_fu_574_p1 = trunc_ln7_reg_733_pp0_iter13_reg;

    assign grp_fu_221_p_ce = 1'b1;

    assign grp_fu_221_p_din0 = grp_fu_274_p0;

    assign grp_fu_221_p_din1 = grp_fu_274_p1;

    assign grp_fu_597_p_ce = 1'b1;

    assign grp_fu_597_p_din0 = grp_fu_257_p0;

    assign grp_fu_597_p_din1 = grp_fu_257_p1;

    assign grp_fu_597_p_opcode = grp_fu_257_opcode;

    assign grp_fu_605_p_ce = 1'b1;

    assign grp_fu_605_p_din0 = grp_fu_262_p0;

    assign grp_fu_605_p_din1 = grp_fu_262_p1;

    assign grp_fu_609_p_ce = 1'b1;

    assign grp_fu_609_p_din0 = grp_fu_267_p0;

    assign grp_fu_609_p_din1 = grp_fu_267_p1;

    assign grp_fu_613_p_ce = 1'b1;

    assign grp_fu_613_p_din0 = laserReading_load_reg_682;

    assign grp_fu_616_p_ce = 1'b1;

    assign grp_fu_616_p_din0 = laserReading_load_reg_682;

    assign grp_fu_616_p_din1 = 32'd0;

    assign grp_fu_616_p_opcode = 5'd3;

    assign grp_fu_620_p_ce = 1'b1;

    assign grp_fu_620_p_din0 = readDist_reg_699;

    assign grp_fu_620_p_din1 = grp_fu_279_p1;

    assign grp_fu_620_p_opcode = grp_fu_279_opcode;

    assign grp_fu_646_p_ce = 1'b1;

    assign grp_fu_646_p_din0 = 64'd0;

    assign grp_fu_646_p_din1 = mul36_i_reg_799_pp0_iter6_reg;

    assign icmp_ln173_fu_311_p2 = ((ap_sig_allocacmp_eIdx_1 == 8'd180) ? 1'b1 : 1'b0);

    assign icmp_ln188_1_fu_387_p2 = ((trunc_ln188_fu_377_p1 == 23'd0) ? 1'b1 : 1'b0);

    assign icmp_ln188_2_fu_429_p2 = ((tmp_7_fu_406_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln188_3_fu_435_p2 = ((trunc_ln188_1_fu_416_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln188_4_fu_447_p2 = ((tmp_8_fu_420_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln188_5_fu_348_p2 = ((trunc_ln188_2 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln188_fu_381_p2 = ((tmp_5_fu_367_p4 != 8'd255) ? 1'b1 : 1'b0);

    assign icmp_ln198_1_fu_498_p2 = ((trunc_ln198_fu_488_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln198_fu_492_p2 = ((tmp_2_fu_478_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign laserReading_address0 = zext_ln177_fu_343_p1;

    assign or_ln188_1_fu_441_p2 = (icmp_ln188_3_fu_435_p2 | icmp_ln188_2_fu_429_p2);

    assign or_ln188_2_fu_453_p2 = (icmp_ln188_5_reg_669 | icmp_ln188_4_fu_447_p2);

    assign or_ln188_fu_393_p2 = (icmp_ln188_reg_689 | icmp_ln188_1_reg_694);

    assign or_ln198_fu_504_p2 = (icmp_ln198_fu_492_p2 | icmp_ln198_1_fu_498_p2);

    assign pMax_fu_566_p3 = ((and_ln193_fu_562_p2[0:0] == 1'b1) ? 64'd4607182418800017408 : 64'd0);

    assign pRand_1_fu_555_p3 = ((and_ln188_fu_550_p2[0:0] == 1'b1) ? pRand : 64'd0);

    assign probability_out = probability_fu_118;

    assign tmp_2_fu_478_p4 = {{bitcast_ln198_fu_475_p1[62:52]}};

    assign tmp_5_fu_367_p4 = {{bitcast_ln188_fu_364_p1[30:23]}};

    assign tmp_7_fu_406_p4 = {{bitcast_ln188_1_fu_403_p1[62:52]}};

    assign tmp_8_fu_420_p4 = {{pf_load_2[254:244]}};

    assign trunc_ln188_1_fu_416_p1 = bitcast_ln188_1_fu_403_p1[51:0];

    assign trunc_ln188_fu_377_p1 = bitcast_ln188_fu_364_p1[22:0];

    assign trunc_ln198_fu_488_p1 = bitcast_ln198_fu_475_p1[51:0];

    assign trunc_ln7_fu_526_p4 = {{pf_load_2[127:64]}};

    assign xor_ln199_fu_535_p2 = (trunc_ln7_fu_526_p4 ^ 64'd9223372036854775808);

    assign zStar_address0 = zext_ln173_fu_326_p1;

    assign zext_ln173_fu_326_p1 = ap_sig_allocacmp_eIdx_1;

    assign zext_ln177_fu_343_p1 = add_ln177_fu_337_p2;

    always @(posedge ap_clk) begin
        pMax_reg_758[51:0]  <= 52'b0000000000000000000000000000000000000000000000000000;
        pMax_reg_758[63:62] <= 2'b00;
    end

endmodule  //main_updateSensor_Pipeline_VITIS_LOOP_173_3
