/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_46_1_VITIS_LOOP_47_2 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    ogm_grid_address0,
    ogm_grid_ce0,
    ogm_grid_we0,
    ogm_grid_d0
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [13:0] ogm_grid_address0;
    output ogm_grid_ce0;
    output ogm_grid_we0;
    output [63:0] ogm_grid_d0;

    reg ap_idle;
    reg ogm_grid_ce0;
    reg ogm_grid_we0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln46_fu_82_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    wire   [6:0] select_ln46_fu_112_p3;
    reg   [6:0] select_ln46_reg_194;
    reg   [6:0] select_ln46_reg_194_pp0_iter1_reg;
    wire   [63:0] zext_ln48_2_fu_156_p1;
    wire    ap_block_pp0_stage0;
    reg   [6:0] j_fu_38;
    wire   [6:0] add_ln47_fu_132_p2;
    wire    ap_loop_init;
    reg   [6:0] ap_sig_allocacmp_j_load;
    reg   [6:0] i_fu_42;
    wire   [6:0] select_ln46_1_fu_120_p3;
    reg   [6:0] ap_sig_allocacmp_i_load;
    reg   [13:0] indvar_flatten_fu_46;
    wire   [13:0] add_ln46_1_fu_88_p2;
    reg   [13:0] ap_sig_allocacmp_indvar_flatten_load;
    wire   [0:0] icmp_ln47_fu_106_p2;
    wire   [6:0] add_ln46_fu_100_p2;
    wire   [13:0] grp_fu_160_p3;
    wire   [6:0] grp_fu_160_p0;
    wire   [6:0] grp_fu_160_p1;
    wire   [6:0] grp_fu_160_p2;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire   [13:0] grp_fu_160_p00;
    wire   [13:0] grp_fu_160_p20;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 j_fu_38 = 7'd0;
        #0 i_fu_42 = 7'd0;
        #0 indvar_flatten_fu_46 = 14'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_mac_muladd_7ns_7ns_7ns_14_4_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(7),
        .din1_WIDTH(7),
        .din2_WIDTH(7),
        .dout_WIDTH(14)
    ) mac_muladd_7ns_7ns_7ns_14_4_1_U1 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_160_p0),
        .din1(grp_fu_160_p1),
        .din2(grp_fu_160_p2),
        .ce(1'b1),
        .dout(grp_fu_160_p3)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln46_fu_82_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                i_fu_42 <= select_ln46_1_fu_120_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                i_fu_42 <= 7'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln46_fu_82_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                indvar_flatten_fu_46 <= add_ln46_1_fu_88_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                indvar_flatten_fu_46 <= 14'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln46_fu_82_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                j_fu_38 <= add_ln47_fu_132_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                j_fu_38 <= 7'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
            select_ln46_reg_194 <= select_ln46_fu_112_p3;
            select_ln46_reg_194_pp0_iter1_reg <= select_ln46_reg_194;
        end
    end

    always @(*) begin
        if (((icmp_ln46_fu_82_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_i_load = 7'd0;
        end else begin
            ap_sig_allocacmp_i_load = i_fu_42;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_indvar_flatten_load = 14'd0;
        end else begin
            ap_sig_allocacmp_indvar_flatten_load = indvar_flatten_fu_46;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_j_load = 7'd0;
        end else begin
            ap_sig_allocacmp_j_load = j_fu_38;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
            ogm_grid_ce0 = 1'b1;
        end else begin
            ogm_grid_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
            ogm_grid_we0 = 1'b1;
        end else begin
            ogm_grid_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln46_1_fu_88_p2 = (ap_sig_allocacmp_indvar_flatten_load + 14'd1);

    assign add_ln46_fu_100_p2 = (ap_sig_allocacmp_i_load + 7'd1);

    assign add_ln47_fu_132_p2 = (select_ln46_fu_112_p3 + 7'd1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign grp_fu_160_p0 = grp_fu_160_p00;

    assign grp_fu_160_p00 = select_ln46_1_fu_120_p3;

    assign grp_fu_160_p1 = 14'd100;

    assign grp_fu_160_p2 = grp_fu_160_p20;

    assign grp_fu_160_p20 = select_ln46_reg_194_pp0_iter1_reg;

    assign icmp_ln46_fu_82_p2 = ((ap_sig_allocacmp_indvar_flatten_load == 14'd10000) ? 1'b1 : 1'b0);

    assign icmp_ln47_fu_106_p2 = ((ap_sig_allocacmp_j_load == 7'd100) ? 1'b1 : 1'b0);

    assign ogm_grid_address0 = zext_ln48_2_fu_156_p1;

    assign ogm_grid_d0 = 64'd4602678819172646912;

    assign select_ln46_1_fu_120_p3 = ((icmp_ln47_fu_106_p2[0:0] == 1'b1) ? add_ln46_fu_100_p2 : ap_sig_allocacmp_i_load);

    assign select_ln46_fu_112_p3 = ((icmp_ln47_fu_106_p2[0:0] == 1'b1) ? 7'd0 : ap_sig_allocacmp_j_load);

    assign zext_ln48_2_fu_156_p1 = grp_fu_160_p3;

endmodule  //main_main_Pipeline_VITIS_LOOP_46_1_VITIS_LOOP_47_2
