/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_detectCollNode (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    this_env_0_0_0_address0,
    this_env_0_0_0_ce0,
    this_env_0_0_0_q0,
    this_env_0_0_1_address0,
    this_env_0_0_1_ce0,
    this_env_0_0_1_q0,
    this_env_0_0_2_address0,
    this_env_0_0_2_ce0,
    this_env_0_0_2_q0,
    this_env_0_1_0_address0,
    this_env_0_1_0_ce0,
    this_env_0_1_0_q0,
    this_env_0_1_1_address0,
    this_env_0_1_1_ce0,
    this_env_0_1_1_q0,
    this_env_0_1_2_address0,
    this_env_0_1_2_ce0,
    this_env_0_1_2_q0,
    this_env_0_2_0_address0,
    this_env_0_2_0_ce0,
    this_env_0_2_0_q0,
    this_env_0_2_1_address0,
    this_env_0_2_1_ce0,
    this_env_0_2_1_q0,
    this_env_0_2_2_address0,
    this_env_0_2_2_ce0,
    this_env_0_2_2_q0,
    this_env_0_3_0_address0,
    this_env_0_3_0_ce0,
    this_env_0_3_0_q0,
    this_env_0_3_1_address0,
    this_env_0_3_1_ce0,
    this_env_0_3_1_q0,
    this_env_0_3_2_address0,
    this_env_0_3_2_ce0,
    this_env_0_3_2_q0,
    this_env_0_4_0_address0,
    this_env_0_4_0_ce0,
    this_env_0_4_0_q0,
    this_env_0_4_1_address0,
    this_env_0_4_1_ce0,
    this_env_0_4_1_q0,
    this_env_0_4_2_address0,
    this_env_0_4_2_ce0,
    this_env_0_4_2_q0,
    this_env_0_5_0_address0,
    this_env_0_5_0_ce0,
    this_env_0_5_0_q0,
    this_env_0_5_1_address0,
    this_env_0_5_1_ce0,
    this_env_0_5_1_q0,
    this_env_0_5_2_address0,
    this_env_0_5_2_ce0,
    this_env_0_5_2_q0,
    this_env_0_6_0_address0,
    this_env_0_6_0_ce0,
    this_env_0_6_0_q0,
    this_env_0_6_1_address0,
    this_env_0_6_1_ce0,
    this_env_0_6_1_q0,
    this_env_0_6_2_address0,
    this_env_0_6_2_ce0,
    this_env_0_6_2_q0,
    this_env_0_7_0_address0,
    this_env_0_7_0_ce0,
    this_env_0_7_0_q0,
    this_env_0_7_1_address0,
    this_env_0_7_1_ce0,
    this_env_0_7_1_q0,
    this_env_0_7_2_address0,
    this_env_0_7_2_ce0,
    this_env_0_7_2_q0,
    this_env_0_8_0_address0,
    this_env_0_8_0_ce0,
    this_env_0_8_0_q0,
    this_env_0_8_1_address0,
    this_env_0_8_1_ce0,
    this_env_0_8_1_q0,
    this_env_0_8_2_address0,
    this_env_0_8_2_ce0,
    this_env_0_8_2_q0,
    this_env_1_address0,
    this_env_1_ce0,
    this_env_1_q0,
    this_env_1_address1,
    this_env_1_ce1,
    this_env_1_q1,
    this_TLink_0_0_address0,
    this_TLink_0_0_ce0,
    this_TLink_0_0_q0,
    this_TLink_0_1_address0,
    this_TLink_0_1_ce0,
    this_TLink_0_1_q0,
    this_TLink_0_2_address0,
    this_TLink_0_2_ce0,
    this_TLink_0_2_q0,
    this_TLink_0_3_address0,
    this_TLink_0_3_ce0,
    this_TLink_0_3_q0,
    this_TLink_1_0_address0,
    this_TLink_1_0_ce0,
    this_TLink_1_0_q0,
    this_TLink_1_1_address0,
    this_TLink_1_1_ce0,
    this_TLink_1_1_q0,
    this_TLink_1_2_address0,
    this_TLink_1_2_ce0,
    this_TLink_1_2_q0,
    this_TLink_1_3_address0,
    this_TLink_1_3_ce0,
    this_TLink_1_3_q0,
    this_TLink_2_0_address0,
    this_TLink_2_0_ce0,
    this_TLink_2_0_q0,
    this_TLink_2_1_address0,
    this_TLink_2_1_ce0,
    this_TLink_2_1_q0,
    this_TLink_2_2_address0,
    this_TLink_2_2_ce0,
    this_TLink_2_2_q0,
    this_TLink_2_3_address0,
    this_TLink_2_3_ce0,
    this_TLink_2_3_q0,
    this_TLink_3_0_address0,
    this_TLink_3_0_ce0,
    this_TLink_3_0_q0,
    this_TLink_3_1_address0,
    this_TLink_3_1_ce0,
    this_TLink_3_1_q0,
    this_TLink_3_2_address0,
    this_TLink_3_2_ce0,
    this_TLink_3_2_q0,
    this_TLink_3_3_address0,
    this_TLink_3_3_ce0,
    this_TLink_3_3_q0,
    this_TJoint_0_0_address0,
    this_TJoint_0_0_ce0,
    this_TJoint_0_0_we0,
    this_TJoint_0_0_d0,
    this_TJoint_0_0_q0,
    this_TJoint_0_1_address0,
    this_TJoint_0_1_ce0,
    this_TJoint_0_1_we0,
    this_TJoint_0_1_d0,
    this_TJoint_0_1_q0,
    this_TJoint_0_2_address0,
    this_TJoint_0_2_ce0,
    this_TJoint_0_2_we0,
    this_TJoint_0_2_d0,
    this_TJoint_0_2_q0,
    this_TJoint_0_3_address0,
    this_TJoint_0_3_ce0,
    this_TJoint_0_3_we0,
    this_TJoint_0_3_d0,
    this_TJoint_0_3_q0,
    this_TJoint_1_0_address0,
    this_TJoint_1_0_ce0,
    this_TJoint_1_0_we0,
    this_TJoint_1_0_d0,
    this_TJoint_1_0_q0,
    this_TJoint_1_1_address0,
    this_TJoint_1_1_ce0,
    this_TJoint_1_1_we0,
    this_TJoint_1_1_d0,
    this_TJoint_1_1_q0,
    this_TJoint_1_2_address0,
    this_TJoint_1_2_ce0,
    this_TJoint_1_2_we0,
    this_TJoint_1_2_d0,
    this_TJoint_1_2_q0,
    this_TJoint_1_3_address0,
    this_TJoint_1_3_ce0,
    this_TJoint_1_3_we0,
    this_TJoint_1_3_d0,
    this_TJoint_1_3_q0,
    this_TJoint_2_0_address0,
    this_TJoint_2_0_ce0,
    this_TJoint_2_0_we0,
    this_TJoint_2_0_d0,
    this_TJoint_2_0_q0,
    this_TJoint_2_1_address0,
    this_TJoint_2_1_ce0,
    this_TJoint_2_1_we0,
    this_TJoint_2_1_d0,
    this_TJoint_2_1_q0,
    this_TJoint_2_2_address0,
    this_TJoint_2_2_ce0,
    this_TJoint_2_2_we0,
    this_TJoint_2_2_d0,
    this_TJoint_2_2_q0,
    this_TJoint_2_3_address0,
    this_TJoint_2_3_ce0,
    this_TJoint_2_3_we0,
    this_TJoint_2_3_d0,
    this_TJoint_2_3_q0,
    this_TJoint_3_0_address0,
    this_TJoint_3_0_ce0,
    this_TJoint_3_0_we0,
    this_TJoint_3_0_d0,
    this_TJoint_3_0_q0,
    this_TJoint_3_1_address0,
    this_TJoint_3_1_ce0,
    this_TJoint_3_1_we0,
    this_TJoint_3_1_d0,
    this_TJoint_3_1_q0,
    this_TJoint_3_2_address0,
    this_TJoint_3_2_ce0,
    this_TJoint_3_2_we0,
    this_TJoint_3_2_d0,
    this_TJoint_3_2_q0,
    this_TJoint_3_3_address0,
    this_TJoint_3_3_ce0,
    this_TJoint_3_3_we0,
    this_TJoint_3_3_d0,
    this_TJoint_3_3_q0,
    this_TCurr_0_0_address0,
    this_TCurr_0_0_ce0,
    this_TCurr_0_0_we0,
    this_TCurr_0_0_d0,
    this_TCurr_0_0_q0,
    this_TCurr_0_1_address0,
    this_TCurr_0_1_ce0,
    this_TCurr_0_1_we0,
    this_TCurr_0_1_d0,
    this_TCurr_0_1_q0,
    this_TCurr_0_2_address0,
    this_TCurr_0_2_ce0,
    this_TCurr_0_2_we0,
    this_TCurr_0_2_d0,
    this_TCurr_0_2_q0,
    this_TCurr_0_3_address0,
    this_TCurr_0_3_ce0,
    this_TCurr_0_3_we0,
    this_TCurr_0_3_d0,
    this_TCurr_0_3_q0,
    this_TCurr_1_0_address0,
    this_TCurr_1_0_ce0,
    this_TCurr_1_0_we0,
    this_TCurr_1_0_d0,
    this_TCurr_1_0_q0,
    this_TCurr_1_1_address0,
    this_TCurr_1_1_ce0,
    this_TCurr_1_1_we0,
    this_TCurr_1_1_d0,
    this_TCurr_1_1_q0,
    this_TCurr_1_2_address0,
    this_TCurr_1_2_ce0,
    this_TCurr_1_2_we0,
    this_TCurr_1_2_d0,
    this_TCurr_1_2_q0,
    this_TCurr_1_3_address0,
    this_TCurr_1_3_ce0,
    this_TCurr_1_3_we0,
    this_TCurr_1_3_d0,
    this_TCurr_1_3_q0,
    this_TCurr_2_0_address0,
    this_TCurr_2_0_ce0,
    this_TCurr_2_0_we0,
    this_TCurr_2_0_d0,
    this_TCurr_2_0_q0,
    this_TCurr_2_1_address0,
    this_TCurr_2_1_ce0,
    this_TCurr_2_1_we0,
    this_TCurr_2_1_d0,
    this_TCurr_2_1_q0,
    this_TCurr_2_2_address0,
    this_TCurr_2_2_ce0,
    this_TCurr_2_2_we0,
    this_TCurr_2_2_d0,
    this_TCurr_2_2_q0,
    this_TCurr_2_3_address0,
    this_TCurr_2_3_ce0,
    this_TCurr_2_3_we0,
    this_TCurr_2_3_d0,
    this_TCurr_2_3_q0,
    this_TCurr_3_0_address0,
    this_TCurr_3_0_ce0,
    this_TCurr_3_0_we0,
    this_TCurr_3_0_d0,
    this_TCurr_3_0_q0,
    this_TCurr_3_1_address0,
    this_TCurr_3_1_ce0,
    this_TCurr_3_1_we0,
    this_TCurr_3_1_d0,
    this_TCurr_3_1_q0,
    this_TCurr_3_2_address0,
    this_TCurr_3_2_ce0,
    this_TCurr_3_2_we0,
    this_TCurr_3_2_d0,
    this_TCurr_3_2_q0,
    this_TCurr_3_3_address0,
    this_TCurr_3_3_ce0,
    this_TCurr_3_3_we0,
    this_TCurr_3_3_d0,
    this_TCurr_3_3_q0,
    this_q_address0,
    this_q_ce0,
    this_q_we0,
    this_q_d0,
    this_q_q0,
    p_read,
    p_read1,
    p_read2,
    p_read3,
    p_read4,
    p_read5,
    p_read6,
    p_read7,
    p_read8,
    p_read9,
    p_read10,
    p_read11,
    p_read12,
    p_read13,
    p_read14,
    p_read15,
    p_read16,
    p_read17,
    p_read18,
    p_read19,
    p_read20,
    p_read21,
    p_read22,
    p_read23,
    p_read24,
    p_read25,
    p_read26,
    p_read27,
    p_read28,
    p_read29,
    p_read30,
    p_read31,
    p_read32,
    p_read33,
    p_read34,
    p_read35,
    p_read36,
    p_read37,
    p_read38,
    p_read39,
    p_read40,
    p_read41,
    p_read42,
    p_read43,
    p_read44,
    p_read45,
    p_read46,
    p_read47,
    p_read48,
    p_read49,
    p_read50,
    p_read51,
    p_read52,
    p_read53,
    p_read54,
    p_read55,
    p_read56,
    p_read57,
    p_read58,
    p_read59,
    p_read60,
    p_read61,
    p_read62,
    p_read63,
    this_cPoints_address0,
    this_cPoints_ce0,
    this_cPoints_we0,
    this_cPoints_d0,
    this_cPoints_q0,
    this_cPoints_address1,
    this_cPoints_ce1,
    this_cPoints_we1,
    this_cPoints_d1,
    this_cPoints_q1,
    this_cAxes_address0,
    this_cAxes_ce0,
    this_cAxes_we0,
    this_cAxes_d0,
    this_cAxes_q0,
    this_cAxes_address1,
    this_cAxes_ce1,
    this_cAxes_q1,
    ang_address0,
    ang_ce0,
    ang_q0,
    l_TColl_0_0_0_constprop_i,
    l_TColl_0_0_0_constprop_o,
    l_TColl_0_0_0_constprop_o_ap_vld,
    l_TColl_0_0_1_constprop_i,
    l_TColl_0_0_1_constprop_o,
    l_TColl_0_0_1_constprop_o_ap_vld,
    l_TColl_0_0_2_constprop_i,
    l_TColl_0_0_2_constprop_o,
    l_TColl_0_0_2_constprop_o_ap_vld,
    l_TColl_0_0_3_constprop_i,
    l_TColl_0_0_3_constprop_o,
    l_TColl_0_0_3_constprop_o_ap_vld,
    l_TColl_1_0_0_constprop_i,
    l_TColl_1_0_0_constprop_o,
    l_TColl_1_0_0_constprop_o_ap_vld,
    l_TColl_1_0_1_constprop_i,
    l_TColl_1_0_1_constprop_o,
    l_TColl_1_0_1_constprop_o_ap_vld,
    l_TColl_1_0_2_constprop_i,
    l_TColl_1_0_2_constprop_o,
    l_TColl_1_0_2_constprop_o_ap_vld,
    l_TColl_1_0_3_constprop_i,
    l_TColl_1_0_3_constprop_o,
    l_TColl_1_0_3_constprop_o_ap_vld,
    l_TColl_2_0_0_constprop_i,
    l_TColl_2_0_0_constprop_o,
    l_TColl_2_0_0_constprop_o_ap_vld,
    l_TColl_2_0_1_constprop_i,
    l_TColl_2_0_1_constprop_o,
    l_TColl_2_0_1_constprop_o_ap_vld,
    l_TColl_2_0_2_constprop_i,
    l_TColl_2_0_2_constprop_o,
    l_TColl_2_0_2_constprop_o_ap_vld,
    l_TColl_2_0_3_constprop_i,
    l_TColl_2_0_3_constprop_o,
    l_TColl_2_0_3_constprop_o_ap_vld,
    l_TColl_0_1_0_constprop_i,
    l_TColl_0_1_0_constprop_o,
    l_TColl_0_1_0_constprop_o_ap_vld,
    l_TColl_0_1_1_constprop_i,
    l_TColl_0_1_1_constprop_o,
    l_TColl_0_1_1_constprop_o_ap_vld,
    l_TColl_0_1_2_constprop_i,
    l_TColl_0_1_2_constprop_o,
    l_TColl_0_1_2_constprop_o_ap_vld,
    l_TColl_0_1_3_constprop_i,
    l_TColl_0_1_3_constprop_o,
    l_TColl_0_1_3_constprop_o_ap_vld,
    l_TColl_1_1_0_constprop_i,
    l_TColl_1_1_0_constprop_o,
    l_TColl_1_1_0_constprop_o_ap_vld,
    l_TColl_1_1_1_constprop_i,
    l_TColl_1_1_1_constprop_o,
    l_TColl_1_1_1_constprop_o_ap_vld,
    l_TColl_1_1_2_constprop_i,
    l_TColl_1_1_2_constprop_o,
    l_TColl_1_1_2_constprop_o_ap_vld,
    l_TColl_1_1_3_constprop_i,
    l_TColl_1_1_3_constprop_o,
    l_TColl_1_1_3_constprop_o_ap_vld,
    l_TColl_2_1_0_constprop_i,
    l_TColl_2_1_0_constprop_o,
    l_TColl_2_1_0_constprop_o_ap_vld,
    l_TColl_2_1_1_constprop_i,
    l_TColl_2_1_1_constprop_o,
    l_TColl_2_1_1_constprop_o_ap_vld,
    l_TColl_2_1_2_constprop_i,
    l_TColl_2_1_2_constprop_o,
    l_TColl_2_1_2_constprop_o_ap_vld,
    l_TColl_2_1_3_constprop_i,
    l_TColl_2_1_3_constprop_o,
    l_TColl_2_1_3_constprop_o_ap_vld,
    l_TColl_0_2_0_constprop_i,
    l_TColl_0_2_0_constprop_o,
    l_TColl_0_2_0_constprop_o_ap_vld,
    l_TColl_0_2_1_constprop_i,
    l_TColl_0_2_1_constprop_o,
    l_TColl_0_2_1_constprop_o_ap_vld,
    l_TColl_0_2_2_constprop_i,
    l_TColl_0_2_2_constprop_o,
    l_TColl_0_2_2_constprop_o_ap_vld,
    l_TColl_0_2_3_constprop_i,
    l_TColl_0_2_3_constprop_o,
    l_TColl_0_2_3_constprop_o_ap_vld,
    l_TColl_1_2_0_constprop_i,
    l_TColl_1_2_0_constprop_o,
    l_TColl_1_2_0_constprop_o_ap_vld,
    l_TColl_1_2_1_constprop_i,
    l_TColl_1_2_1_constprop_o,
    l_TColl_1_2_1_constprop_o_ap_vld,
    l_TColl_1_2_2_constprop_i,
    l_TColl_1_2_2_constprop_o,
    l_TColl_1_2_2_constprop_o_ap_vld,
    l_TColl_1_2_3_constprop_i,
    l_TColl_1_2_3_constprop_o,
    l_TColl_1_2_3_constprop_o_ap_vld,
    l_TColl_2_2_0_constprop_i,
    l_TColl_2_2_0_constprop_o,
    l_TColl_2_2_0_constprop_o_ap_vld,
    l_TColl_2_2_1_constprop_i,
    l_TColl_2_2_1_constprop_o,
    l_TColl_2_2_1_constprop_o_ap_vld,
    l_TColl_2_2_2_constprop_i,
    l_TColl_2_2_2_constprop_o,
    l_TColl_2_2_2_constprop_o_ap_vld,
    l_TColl_2_2_3_constprop_i,
    l_TColl_2_2_3_constprop_o,
    l_TColl_2_2_3_constprop_o_ap_vld,
    l_TColl_0_3_0_constprop_i,
    l_TColl_0_3_0_constprop_o,
    l_TColl_0_3_0_constprop_o_ap_vld,
    l_TColl_0_3_1_constprop_i,
    l_TColl_0_3_1_constprop_o,
    l_TColl_0_3_1_constprop_o_ap_vld,
    l_TColl_0_3_2_constprop_i,
    l_TColl_0_3_2_constprop_o,
    l_TColl_0_3_2_constprop_o_ap_vld,
    l_TColl_0_3_3_constprop_i,
    l_TColl_0_3_3_constprop_o,
    l_TColl_0_3_3_constprop_o_ap_vld,
    l_TColl_1_3_0_constprop_i,
    l_TColl_1_3_0_constprop_o,
    l_TColl_1_3_0_constprop_o_ap_vld,
    l_TColl_1_3_1_constprop_i,
    l_TColl_1_3_1_constprop_o,
    l_TColl_1_3_1_constprop_o_ap_vld,
    l_TColl_1_3_2_constprop_i,
    l_TColl_1_3_2_constprop_o,
    l_TColl_1_3_2_constprop_o_ap_vld,
    l_TColl_1_3_3_constprop_i,
    l_TColl_1_3_3_constprop_o,
    l_TColl_1_3_3_constprop_o_ap_vld,
    l_TColl_2_3_0_constprop_i,
    l_TColl_2_3_0_constprop_o,
    l_TColl_2_3_0_constprop_o_ap_vld,
    l_TColl_2_3_1_constprop_i,
    l_TColl_2_3_1_constprop_o,
    l_TColl_2_3_1_constprop_o_ap_vld,
    l_TColl_2_3_2_constprop_i,
    l_TColl_2_3_2_constprop_o,
    l_TColl_2_3_2_constprop_o_ap_vld,
    l_TColl_2_3_3_constprop_i,
    l_TColl_2_3_3_constprop_o,
    l_TColl_2_3_3_constprop_o_ap_vld,
    ap_return,
    grp_fu_2529_p_din0,
    grp_fu_2529_p_din1,
    grp_fu_2529_p_opcode,
    grp_fu_2529_p_dout0,
    grp_fu_2529_p_ce,
    grp_fu_2533_p_din0,
    grp_fu_2533_p_din1,
    grp_fu_2533_p_dout0,
    grp_fu_2533_p_ce,
    grp_fu_2537_p_din0,
    grp_fu_2537_p_din1,
    grp_fu_2537_p_opcode,
    grp_fu_2537_p_dout0,
    grp_fu_2537_p_ce,
    grp_fu_2541_p_din0,
    grp_fu_2541_p_din1,
    grp_fu_2541_p_opcode,
    grp_fu_2541_p_dout0,
    grp_fu_2541_p_ce,
    grp_fu_2545_p_din0,
    grp_fu_2545_p_din1,
    grp_fu_2545_p_opcode,
    grp_fu_2545_p_dout0,
    grp_fu_2545_p_ce,
    grp_fu_2549_p_din0,
    grp_fu_2549_p_din1,
    grp_fu_2549_p_opcode,
    grp_fu_2549_p_dout0,
    grp_fu_2549_p_ce,
    grp_fu_2553_p_din0,
    grp_fu_2553_p_din1,
    grp_fu_2553_p_opcode,
    grp_fu_2553_p_dout0,
    grp_fu_2553_p_ce,
    grp_fu_2557_p_din0,
    grp_fu_2557_p_din1,
    grp_fu_2557_p_dout0,
    grp_fu_2557_p_ce,
    grp_fu_2561_p_din0,
    grp_fu_2561_p_din1,
    grp_fu_2561_p_dout0,
    grp_fu_2561_p_ce,
    grp_fu_2565_p_din0,
    grp_fu_2565_p_din1,
    grp_fu_2565_p_dout0,
    grp_fu_2565_p_ce,
    grp_fu_1454_p_din0,
    grp_fu_1454_p_din1,
    grp_fu_1454_p_opcode,
    grp_fu_1454_p_dout0,
    grp_fu_1454_p_ce,
    grp_fu_1462_p_din0,
    grp_fu_1462_p_din1,
    grp_fu_1462_p_dout0,
    grp_fu_1462_p_ce
);

    parameter ap_ST_fsm_state1 = 8'd1;
    parameter ap_ST_fsm_state2 = 8'd2;
    parameter ap_ST_fsm_state3 = 8'd4;
    parameter ap_ST_fsm_state4 = 8'd8;
    parameter ap_ST_fsm_state5 = 8'd16;
    parameter ap_ST_fsm_state6 = 8'd32;
    parameter ap_ST_fsm_state7 = 8'd64;
    parameter ap_ST_fsm_state8 = 8'd128;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [2:0] this_env_0_0_0_address0;
    output this_env_0_0_0_ce0;
    input [63:0] this_env_0_0_0_q0;
    output [2:0] this_env_0_0_1_address0;
    output this_env_0_0_1_ce0;
    input [63:0] this_env_0_0_1_q0;
    output [2:0] this_env_0_0_2_address0;
    output this_env_0_0_2_ce0;
    input [63:0] this_env_0_0_2_q0;
    output [2:0] this_env_0_1_0_address0;
    output this_env_0_1_0_ce0;
    input [63:0] this_env_0_1_0_q0;
    output [2:0] this_env_0_1_1_address0;
    output this_env_0_1_1_ce0;
    input [63:0] this_env_0_1_1_q0;
    output [2:0] this_env_0_1_2_address0;
    output this_env_0_1_2_ce0;
    input [63:0] this_env_0_1_2_q0;
    output [2:0] this_env_0_2_0_address0;
    output this_env_0_2_0_ce0;
    input [63:0] this_env_0_2_0_q0;
    output [2:0] this_env_0_2_1_address0;
    output this_env_0_2_1_ce0;
    input [63:0] this_env_0_2_1_q0;
    output [2:0] this_env_0_2_2_address0;
    output this_env_0_2_2_ce0;
    input [63:0] this_env_0_2_2_q0;
    output [2:0] this_env_0_3_0_address0;
    output this_env_0_3_0_ce0;
    input [63:0] this_env_0_3_0_q0;
    output [2:0] this_env_0_3_1_address0;
    output this_env_0_3_1_ce0;
    input [63:0] this_env_0_3_1_q0;
    output [2:0] this_env_0_3_2_address0;
    output this_env_0_3_2_ce0;
    input [63:0] this_env_0_3_2_q0;
    output [2:0] this_env_0_4_0_address0;
    output this_env_0_4_0_ce0;
    input [63:0] this_env_0_4_0_q0;
    output [2:0] this_env_0_4_1_address0;
    output this_env_0_4_1_ce0;
    input [63:0] this_env_0_4_1_q0;
    output [2:0] this_env_0_4_2_address0;
    output this_env_0_4_2_ce0;
    input [63:0] this_env_0_4_2_q0;
    output [2:0] this_env_0_5_0_address0;
    output this_env_0_5_0_ce0;
    input [63:0] this_env_0_5_0_q0;
    output [2:0] this_env_0_5_1_address0;
    output this_env_0_5_1_ce0;
    input [63:0] this_env_0_5_1_q0;
    output [2:0] this_env_0_5_2_address0;
    output this_env_0_5_2_ce0;
    input [63:0] this_env_0_5_2_q0;
    output [2:0] this_env_0_6_0_address0;
    output this_env_0_6_0_ce0;
    input [63:0] this_env_0_6_0_q0;
    output [2:0] this_env_0_6_1_address0;
    output this_env_0_6_1_ce0;
    input [63:0] this_env_0_6_1_q0;
    output [2:0] this_env_0_6_2_address0;
    output this_env_0_6_2_ce0;
    input [63:0] this_env_0_6_2_q0;
    output [2:0] this_env_0_7_0_address0;
    output this_env_0_7_0_ce0;
    input [63:0] this_env_0_7_0_q0;
    output [2:0] this_env_0_7_1_address0;
    output this_env_0_7_1_ce0;
    input [63:0] this_env_0_7_1_q0;
    output [2:0] this_env_0_7_2_address0;
    output this_env_0_7_2_ce0;
    input [63:0] this_env_0_7_2_q0;
    output [2:0] this_env_0_8_0_address0;
    output this_env_0_8_0_ce0;
    input [63:0] this_env_0_8_0_q0;
    output [2:0] this_env_0_8_1_address0;
    output this_env_0_8_1_ce0;
    input [63:0] this_env_0_8_1_q0;
    output [2:0] this_env_0_8_2_address0;
    output this_env_0_8_2_ce0;
    input [63:0] this_env_0_8_2_q0;
    output [6:0] this_env_1_address0;
    output this_env_1_ce0;
    input [63:0] this_env_1_q0;
    output [6:0] this_env_1_address1;
    output this_env_1_ce1;
    input [63:0] this_env_1_q1;
    output [2:0] this_TLink_0_0_address0;
    output this_TLink_0_0_ce0;
    input [63:0] this_TLink_0_0_q0;
    output [2:0] this_TLink_0_1_address0;
    output this_TLink_0_1_ce0;
    input [63:0] this_TLink_0_1_q0;
    output [2:0] this_TLink_0_2_address0;
    output this_TLink_0_2_ce0;
    input [63:0] this_TLink_0_2_q0;
    output [2:0] this_TLink_0_3_address0;
    output this_TLink_0_3_ce0;
    input [63:0] this_TLink_0_3_q0;
    output [2:0] this_TLink_1_0_address0;
    output this_TLink_1_0_ce0;
    input [63:0] this_TLink_1_0_q0;
    output [2:0] this_TLink_1_1_address0;
    output this_TLink_1_1_ce0;
    input [63:0] this_TLink_1_1_q0;
    output [2:0] this_TLink_1_2_address0;
    output this_TLink_1_2_ce0;
    input [63:0] this_TLink_1_2_q0;
    output [2:0] this_TLink_1_3_address0;
    output this_TLink_1_3_ce0;
    input [63:0] this_TLink_1_3_q0;
    output [2:0] this_TLink_2_0_address0;
    output this_TLink_2_0_ce0;
    input [63:0] this_TLink_2_0_q0;
    output [2:0] this_TLink_2_1_address0;
    output this_TLink_2_1_ce0;
    input [63:0] this_TLink_2_1_q0;
    output [2:0] this_TLink_2_2_address0;
    output this_TLink_2_2_ce0;
    input [63:0] this_TLink_2_2_q0;
    output [2:0] this_TLink_2_3_address0;
    output this_TLink_2_3_ce0;
    input [63:0] this_TLink_2_3_q0;
    output [2:0] this_TLink_3_0_address0;
    output this_TLink_3_0_ce0;
    input [63:0] this_TLink_3_0_q0;
    output [2:0] this_TLink_3_1_address0;
    output this_TLink_3_1_ce0;
    input [63:0] this_TLink_3_1_q0;
    output [2:0] this_TLink_3_2_address0;
    output this_TLink_3_2_ce0;
    input [63:0] this_TLink_3_2_q0;
    output [2:0] this_TLink_3_3_address0;
    output this_TLink_3_3_ce0;
    input [63:0] this_TLink_3_3_q0;
    output [2:0] this_TJoint_0_0_address0;
    output this_TJoint_0_0_ce0;
    output this_TJoint_0_0_we0;
    output [63:0] this_TJoint_0_0_d0;
    input [63:0] this_TJoint_0_0_q0;
    output [2:0] this_TJoint_0_1_address0;
    output this_TJoint_0_1_ce0;
    output this_TJoint_0_1_we0;
    output [63:0] this_TJoint_0_1_d0;
    input [63:0] this_TJoint_0_1_q0;
    output [2:0] this_TJoint_0_2_address0;
    output this_TJoint_0_2_ce0;
    output this_TJoint_0_2_we0;
    output [63:0] this_TJoint_0_2_d0;
    input [63:0] this_TJoint_0_2_q0;
    output [2:0] this_TJoint_0_3_address0;
    output this_TJoint_0_3_ce0;
    output this_TJoint_0_3_we0;
    output [63:0] this_TJoint_0_3_d0;
    input [63:0] this_TJoint_0_3_q0;
    output [2:0] this_TJoint_1_0_address0;
    output this_TJoint_1_0_ce0;
    output this_TJoint_1_0_we0;
    output [63:0] this_TJoint_1_0_d0;
    input [63:0] this_TJoint_1_0_q0;
    output [2:0] this_TJoint_1_1_address0;
    output this_TJoint_1_1_ce0;
    output this_TJoint_1_1_we0;
    output [63:0] this_TJoint_1_1_d0;
    input [63:0] this_TJoint_1_1_q0;
    output [2:0] this_TJoint_1_2_address0;
    output this_TJoint_1_2_ce0;
    output this_TJoint_1_2_we0;
    output [63:0] this_TJoint_1_2_d0;
    input [63:0] this_TJoint_1_2_q0;
    output [2:0] this_TJoint_1_3_address0;
    output this_TJoint_1_3_ce0;
    output this_TJoint_1_3_we0;
    output [63:0] this_TJoint_1_3_d0;
    input [63:0] this_TJoint_1_3_q0;
    output [2:0] this_TJoint_2_0_address0;
    output this_TJoint_2_0_ce0;
    output this_TJoint_2_0_we0;
    output [63:0] this_TJoint_2_0_d0;
    input [63:0] this_TJoint_2_0_q0;
    output [2:0] this_TJoint_2_1_address0;
    output this_TJoint_2_1_ce0;
    output this_TJoint_2_1_we0;
    output [63:0] this_TJoint_2_1_d0;
    input [63:0] this_TJoint_2_1_q0;
    output [2:0] this_TJoint_2_2_address0;
    output this_TJoint_2_2_ce0;
    output this_TJoint_2_2_we0;
    output [63:0] this_TJoint_2_2_d0;
    input [63:0] this_TJoint_2_2_q0;
    output [2:0] this_TJoint_2_3_address0;
    output this_TJoint_2_3_ce0;
    output this_TJoint_2_3_we0;
    output [63:0] this_TJoint_2_3_d0;
    input [63:0] this_TJoint_2_3_q0;
    output [2:0] this_TJoint_3_0_address0;
    output this_TJoint_3_0_ce0;
    output this_TJoint_3_0_we0;
    output [63:0] this_TJoint_3_0_d0;
    input [63:0] this_TJoint_3_0_q0;
    output [2:0] this_TJoint_3_1_address0;
    output this_TJoint_3_1_ce0;
    output this_TJoint_3_1_we0;
    output [63:0] this_TJoint_3_1_d0;
    input [63:0] this_TJoint_3_1_q0;
    output [2:0] this_TJoint_3_2_address0;
    output this_TJoint_3_2_ce0;
    output this_TJoint_3_2_we0;
    output [63:0] this_TJoint_3_2_d0;
    input [63:0] this_TJoint_3_2_q0;
    output [2:0] this_TJoint_3_3_address0;
    output this_TJoint_3_3_ce0;
    output this_TJoint_3_3_we0;
    output [63:0] this_TJoint_3_3_d0;
    input [63:0] this_TJoint_3_3_q0;
    output [2:0] this_TCurr_0_0_address0;
    output this_TCurr_0_0_ce0;
    output this_TCurr_0_0_we0;
    output [63:0] this_TCurr_0_0_d0;
    input [63:0] this_TCurr_0_0_q0;
    output [2:0] this_TCurr_0_1_address0;
    output this_TCurr_0_1_ce0;
    output this_TCurr_0_1_we0;
    output [63:0] this_TCurr_0_1_d0;
    input [63:0] this_TCurr_0_1_q0;
    output [2:0] this_TCurr_0_2_address0;
    output this_TCurr_0_2_ce0;
    output this_TCurr_0_2_we0;
    output [63:0] this_TCurr_0_2_d0;
    input [63:0] this_TCurr_0_2_q0;
    output [2:0] this_TCurr_0_3_address0;
    output this_TCurr_0_3_ce0;
    output this_TCurr_0_3_we0;
    output [63:0] this_TCurr_0_3_d0;
    input [63:0] this_TCurr_0_3_q0;
    output [2:0] this_TCurr_1_0_address0;
    output this_TCurr_1_0_ce0;
    output this_TCurr_1_0_we0;
    output [63:0] this_TCurr_1_0_d0;
    input [63:0] this_TCurr_1_0_q0;
    output [2:0] this_TCurr_1_1_address0;
    output this_TCurr_1_1_ce0;
    output this_TCurr_1_1_we0;
    output [63:0] this_TCurr_1_1_d0;
    input [63:0] this_TCurr_1_1_q0;
    output [2:0] this_TCurr_1_2_address0;
    output this_TCurr_1_2_ce0;
    output this_TCurr_1_2_we0;
    output [63:0] this_TCurr_1_2_d0;
    input [63:0] this_TCurr_1_2_q0;
    output [2:0] this_TCurr_1_3_address0;
    output this_TCurr_1_3_ce0;
    output this_TCurr_1_3_we0;
    output [63:0] this_TCurr_1_3_d0;
    input [63:0] this_TCurr_1_3_q0;
    output [2:0] this_TCurr_2_0_address0;
    output this_TCurr_2_0_ce0;
    output this_TCurr_2_0_we0;
    output [63:0] this_TCurr_2_0_d0;
    input [63:0] this_TCurr_2_0_q0;
    output [2:0] this_TCurr_2_1_address0;
    output this_TCurr_2_1_ce0;
    output this_TCurr_2_1_we0;
    output [63:0] this_TCurr_2_1_d0;
    input [63:0] this_TCurr_2_1_q0;
    output [2:0] this_TCurr_2_2_address0;
    output this_TCurr_2_2_ce0;
    output this_TCurr_2_2_we0;
    output [63:0] this_TCurr_2_2_d0;
    input [63:0] this_TCurr_2_2_q0;
    output [2:0] this_TCurr_2_3_address0;
    output this_TCurr_2_3_ce0;
    output this_TCurr_2_3_we0;
    output [63:0] this_TCurr_2_3_d0;
    input [63:0] this_TCurr_2_3_q0;
    output [2:0] this_TCurr_3_0_address0;
    output this_TCurr_3_0_ce0;
    output this_TCurr_3_0_we0;
    output [63:0] this_TCurr_3_0_d0;
    input [63:0] this_TCurr_3_0_q0;
    output [2:0] this_TCurr_3_1_address0;
    output this_TCurr_3_1_ce0;
    output this_TCurr_3_1_we0;
    output [63:0] this_TCurr_3_1_d0;
    input [63:0] this_TCurr_3_1_q0;
    output [2:0] this_TCurr_3_2_address0;
    output this_TCurr_3_2_ce0;
    output this_TCurr_3_2_we0;
    output [63:0] this_TCurr_3_2_d0;
    input [63:0] this_TCurr_3_2_q0;
    output [2:0] this_TCurr_3_3_address0;
    output this_TCurr_3_3_ce0;
    output this_TCurr_3_3_we0;
    output [63:0] this_TCurr_3_3_d0;
    input [63:0] this_TCurr_3_3_q0;
    output [2:0] this_q_address0;
    output this_q_ce0;
    output this_q_we0;
    output [63:0] this_q_d0;
    input [63:0] this_q_q0;
    input [63:0] p_read;
    input [63:0] p_read1;
    input [63:0] p_read2;
    input [63:0] p_read3;
    input [63:0] p_read4;
    input [63:0] p_read5;
    input [63:0] p_read6;
    input [63:0] p_read7;
    input [63:0] p_read8;
    input [63:0] p_read9;
    input [63:0] p_read10;
    input [63:0] p_read11;
    input [63:0] p_read12;
    input [63:0] p_read13;
    input [63:0] p_read14;
    input [63:0] p_read15;
    input [63:0] p_read16;
    input [63:0] p_read17;
    input [63:0] p_read18;
    input [63:0] p_read19;
    input [63:0] p_read20;
    input [63:0] p_read21;
    input [63:0] p_read22;
    input [63:0] p_read23;
    input [63:0] p_read24;
    input [63:0] p_read25;
    input [63:0] p_read26;
    input [63:0] p_read27;
    input [63:0] p_read28;
    input [63:0] p_read29;
    input [63:0] p_read30;
    input [63:0] p_read31;
    input [63:0] p_read32;
    input [63:0] p_read33;
    input [63:0] p_read34;
    input [63:0] p_read35;
    input [63:0] p_read36;
    input [63:0] p_read37;
    input [63:0] p_read38;
    input [63:0] p_read39;
    input [63:0] p_read40;
    input [63:0] p_read41;
    input [63:0] p_read42;
    input [63:0] p_read43;
    input [63:0] p_read44;
    input [63:0] p_read45;
    input [63:0] p_read46;
    input [63:0] p_read47;
    input [63:0] p_read48;
    input [63:0] p_read49;
    input [63:0] p_read50;
    input [63:0] p_read51;
    input [63:0] p_read52;
    input [63:0] p_read53;
    input [63:0] p_read54;
    input [63:0] p_read55;
    input [63:0] p_read56;
    input [63:0] p_read57;
    input [63:0] p_read58;
    input [63:0] p_read59;
    input [63:0] p_read60;
    input [63:0] p_read61;
    input [63:0] p_read62;
    input [63:0] p_read63;
    output [6:0] this_cPoints_address0;
    output this_cPoints_ce0;
    output this_cPoints_we0;
    output [63:0] this_cPoints_d0;
    input [63:0] this_cPoints_q0;
    output [6:0] this_cPoints_address1;
    output this_cPoints_ce1;
    output this_cPoints_we1;
    output [63:0] this_cPoints_d1;
    input [63:0] this_cPoints_q1;
    output [5:0] this_cAxes_address0;
    output this_cAxes_ce0;
    output this_cAxes_we0;
    output [63:0] this_cAxes_d0;
    input [63:0] this_cAxes_q0;
    output [5:0] this_cAxes_address1;
    output this_cAxes_ce1;
    input [63:0] this_cAxes_q1;
    output [2:0] ang_address0;
    output ang_ce0;
    input [63:0] ang_q0;
    input [63:0] l_TColl_0_0_0_constprop_i;
    output [63:0] l_TColl_0_0_0_constprop_o;
    output l_TColl_0_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_1_constprop_i;
    output [63:0] l_TColl_0_0_1_constprop_o;
    output l_TColl_0_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_2_constprop_i;
    output [63:0] l_TColl_0_0_2_constprop_o;
    output l_TColl_0_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_3_constprop_i;
    output [63:0] l_TColl_0_0_3_constprop_o;
    output l_TColl_0_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_0_constprop_i;
    output [63:0] l_TColl_1_0_0_constprop_o;
    output l_TColl_1_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_1_constprop_i;
    output [63:0] l_TColl_1_0_1_constprop_o;
    output l_TColl_1_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_2_constprop_i;
    output [63:0] l_TColl_1_0_2_constprop_o;
    output l_TColl_1_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_3_constprop_i;
    output [63:0] l_TColl_1_0_3_constprop_o;
    output l_TColl_1_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_0_constprop_i;
    output [63:0] l_TColl_2_0_0_constprop_o;
    output l_TColl_2_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_1_constprop_i;
    output [63:0] l_TColl_2_0_1_constprop_o;
    output l_TColl_2_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_2_constprop_i;
    output [63:0] l_TColl_2_0_2_constprop_o;
    output l_TColl_2_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_3_constprop_i;
    output [63:0] l_TColl_2_0_3_constprop_o;
    output l_TColl_2_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_0_constprop_i;
    output [63:0] l_TColl_0_1_0_constprop_o;
    output l_TColl_0_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_1_constprop_i;
    output [63:0] l_TColl_0_1_1_constprop_o;
    output l_TColl_0_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_2_constprop_i;
    output [63:0] l_TColl_0_1_2_constprop_o;
    output l_TColl_0_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_3_constprop_i;
    output [63:0] l_TColl_0_1_3_constprop_o;
    output l_TColl_0_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_0_constprop_i;
    output [63:0] l_TColl_1_1_0_constprop_o;
    output l_TColl_1_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_1_constprop_i;
    output [63:0] l_TColl_1_1_1_constprop_o;
    output l_TColl_1_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_2_constprop_i;
    output [63:0] l_TColl_1_1_2_constprop_o;
    output l_TColl_1_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_3_constprop_i;
    output [63:0] l_TColl_1_1_3_constprop_o;
    output l_TColl_1_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_0_constprop_i;
    output [63:0] l_TColl_2_1_0_constprop_o;
    output l_TColl_2_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_1_constprop_i;
    output [63:0] l_TColl_2_1_1_constprop_o;
    output l_TColl_2_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_2_constprop_i;
    output [63:0] l_TColl_2_1_2_constprop_o;
    output l_TColl_2_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_3_constprop_i;
    output [63:0] l_TColl_2_1_3_constprop_o;
    output l_TColl_2_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_0_constprop_i;
    output [63:0] l_TColl_0_2_0_constprop_o;
    output l_TColl_0_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_1_constprop_i;
    output [63:0] l_TColl_0_2_1_constprop_o;
    output l_TColl_0_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_2_constprop_i;
    output [63:0] l_TColl_0_2_2_constprop_o;
    output l_TColl_0_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_3_constprop_i;
    output [63:0] l_TColl_0_2_3_constprop_o;
    output l_TColl_0_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_0_constprop_i;
    output [63:0] l_TColl_1_2_0_constprop_o;
    output l_TColl_1_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_1_constprop_i;
    output [63:0] l_TColl_1_2_1_constprop_o;
    output l_TColl_1_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_2_constprop_i;
    output [63:0] l_TColl_1_2_2_constprop_o;
    output l_TColl_1_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_3_constprop_i;
    output [63:0] l_TColl_1_2_3_constprop_o;
    output l_TColl_1_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_0_constprop_i;
    output [63:0] l_TColl_2_2_0_constprop_o;
    output l_TColl_2_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_1_constprop_i;
    output [63:0] l_TColl_2_2_1_constprop_o;
    output l_TColl_2_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_2_constprop_i;
    output [63:0] l_TColl_2_2_2_constprop_o;
    output l_TColl_2_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_3_constprop_i;
    output [63:0] l_TColl_2_2_3_constprop_o;
    output l_TColl_2_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_0_constprop_i;
    output [63:0] l_TColl_0_3_0_constprop_o;
    output l_TColl_0_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_1_constprop_i;
    output [63:0] l_TColl_0_3_1_constprop_o;
    output l_TColl_0_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_2_constprop_i;
    output [63:0] l_TColl_0_3_2_constprop_o;
    output l_TColl_0_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_3_constprop_i;
    output [63:0] l_TColl_0_3_3_constprop_o;
    output l_TColl_0_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_0_constprop_i;
    output [63:0] l_TColl_1_3_0_constprop_o;
    output l_TColl_1_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_1_constprop_i;
    output [63:0] l_TColl_1_3_1_constprop_o;
    output l_TColl_1_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_2_constprop_i;
    output [63:0] l_TColl_1_3_2_constprop_o;
    output l_TColl_1_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_3_constprop_i;
    output [63:0] l_TColl_1_3_3_constprop_o;
    output l_TColl_1_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_0_constprop_i;
    output [63:0] l_TColl_2_3_0_constprop_o;
    output l_TColl_2_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_1_constprop_i;
    output [63:0] l_TColl_2_3_1_constprop_o;
    output l_TColl_2_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_2_constprop_i;
    output [63:0] l_TColl_2_3_2_constprop_o;
    output l_TColl_2_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_3_constprop_i;
    output [63:0] l_TColl_2_3_3_constprop_o;
    output l_TColl_2_3_3_constprop_o_ap_vld;
    output [0:0] ap_return;
    output [63:0] grp_fu_2529_p_din0;
    output [63:0] grp_fu_2529_p_din1;
    output [1:0] grp_fu_2529_p_opcode;
    input [63:0] grp_fu_2529_p_dout0;
    output grp_fu_2529_p_ce;
    output [63:0] grp_fu_2533_p_din0;
    output [63:0] grp_fu_2533_p_din1;
    input [63:0] grp_fu_2533_p_dout0;
    output grp_fu_2533_p_ce;
    output [63:0] grp_fu_2537_p_din0;
    output [63:0] grp_fu_2537_p_din1;
    output [1:0] grp_fu_2537_p_opcode;
    input [63:0] grp_fu_2537_p_dout0;
    output grp_fu_2537_p_ce;
    output [63:0] grp_fu_2541_p_din0;
    output [63:0] grp_fu_2541_p_din1;
    output [1:0] grp_fu_2541_p_opcode;
    input [63:0] grp_fu_2541_p_dout0;
    output grp_fu_2541_p_ce;
    output [63:0] grp_fu_2545_p_din0;
    output [63:0] grp_fu_2545_p_din1;
    output [1:0] grp_fu_2545_p_opcode;
    input [63:0] grp_fu_2545_p_dout0;
    output grp_fu_2545_p_ce;
    output [63:0] grp_fu_2549_p_din0;
    output [63:0] grp_fu_2549_p_din1;
    output [1:0] grp_fu_2549_p_opcode;
    input [63:0] grp_fu_2549_p_dout0;
    output grp_fu_2549_p_ce;
    output [63:0] grp_fu_2553_p_din0;
    output [63:0] grp_fu_2553_p_din1;
    output [1:0] grp_fu_2553_p_opcode;
    input [63:0] grp_fu_2553_p_dout0;
    output grp_fu_2553_p_ce;
    output [63:0] grp_fu_2557_p_din0;
    output [63:0] grp_fu_2557_p_din1;
    input [63:0] grp_fu_2557_p_dout0;
    output grp_fu_2557_p_ce;
    output [63:0] grp_fu_2561_p_din0;
    output [63:0] grp_fu_2561_p_din1;
    input [63:0] grp_fu_2561_p_dout0;
    output grp_fu_2561_p_ce;
    output [63:0] grp_fu_2565_p_din0;
    output [63:0] grp_fu_2565_p_din1;
    input [63:0] grp_fu_2565_p_dout0;
    output grp_fu_2565_p_ce;
    output [63:0] grp_fu_1454_p_din0;
    output [63:0] grp_fu_1454_p_din1;
    output [4:0] grp_fu_1454_p_opcode;
    input [0:0] grp_fu_1454_p_dout0;
    output grp_fu_1454_p_ce;
    output [63:0] grp_fu_1462_p_din0;
    output [63:0] grp_fu_1462_p_din1;
    input [63:0] grp_fu_1462_p_dout0;
    output grp_fu_1462_p_ce;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg [2:0] this_TCurr_0_0_address0;
    reg this_TCurr_0_0_ce0;
    reg this_TCurr_0_0_we0;
    reg [2:0] this_TCurr_0_1_address0;
    reg this_TCurr_0_1_ce0;
    reg this_TCurr_0_1_we0;
    reg [2:0] this_TCurr_0_2_address0;
    reg this_TCurr_0_2_ce0;
    reg this_TCurr_0_2_we0;
    reg [2:0] this_TCurr_0_3_address0;
    reg this_TCurr_0_3_ce0;
    reg this_TCurr_0_3_we0;
    reg [2:0] this_TCurr_1_0_address0;
    reg this_TCurr_1_0_ce0;
    reg this_TCurr_1_0_we0;
    reg [2:0] this_TCurr_1_1_address0;
    reg this_TCurr_1_1_ce0;
    reg this_TCurr_1_1_we0;
    reg [2:0] this_TCurr_1_2_address0;
    reg this_TCurr_1_2_ce0;
    reg this_TCurr_1_2_we0;
    reg [2:0] this_TCurr_1_3_address0;
    reg this_TCurr_1_3_ce0;
    reg this_TCurr_1_3_we0;
    reg [2:0] this_TCurr_2_0_address0;
    reg this_TCurr_2_0_ce0;
    reg this_TCurr_2_0_we0;
    reg [2:0] this_TCurr_2_1_address0;
    reg this_TCurr_2_1_ce0;
    reg this_TCurr_2_1_we0;
    reg [2:0] this_TCurr_2_2_address0;
    reg this_TCurr_2_2_ce0;
    reg this_TCurr_2_2_we0;
    reg [2:0] this_TCurr_2_3_address0;
    reg this_TCurr_2_3_ce0;
    reg this_TCurr_2_3_we0;
    reg [6:0] this_cPoints_address0;
    reg this_cPoints_ce0;
    reg this_cPoints_we0;
    reg [6:0] this_cPoints_address1;
    reg this_cPoints_ce1;
    reg this_cPoints_we1;
    reg [5:0] this_cAxes_address0;
    reg this_cAxes_ce0;
    reg this_cAxes_we0;
    reg this_cAxes_ce1;
    reg [63:0] l_TColl_0_0_0_constprop_o;
    reg [63:0] l_TColl_0_0_1_constprop_o;
    reg [63:0] l_TColl_0_0_2_constprop_o;
    reg [63:0] l_TColl_0_0_3_constprop_o;
    reg [63:0] l_TColl_1_0_0_constprop_o;
    reg [63:0] l_TColl_1_0_1_constprop_o;
    reg [63:0] l_TColl_1_0_2_constprop_o;
    reg [63:0] l_TColl_1_0_3_constprop_o;
    reg [63:0] l_TColl_2_0_0_constprop_o;
    reg [63:0] l_TColl_2_0_1_constprop_o;
    reg [63:0] l_TColl_2_0_2_constprop_o;
    reg [63:0] l_TColl_2_0_3_constprop_o;
    reg [63:0] l_TColl_0_1_0_constprop_o;
    reg [63:0] l_TColl_0_1_1_constprop_o;
    reg [63:0] l_TColl_0_1_2_constprop_o;
    reg [63:0] l_TColl_0_1_3_constprop_o;
    reg [63:0] l_TColl_1_1_0_constprop_o;
    reg [63:0] l_TColl_1_1_1_constprop_o;
    reg [63:0] l_TColl_1_1_2_constprop_o;
    reg [63:0] l_TColl_1_1_3_constprop_o;
    reg [63:0] l_TColl_2_1_0_constprop_o;
    reg [63:0] l_TColl_2_1_1_constprop_o;
    reg [63:0] l_TColl_2_1_2_constprop_o;
    reg [63:0] l_TColl_2_1_3_constprop_o;
    reg [63:0] l_TColl_0_2_0_constprop_o;
    reg [63:0] l_TColl_0_2_1_constprop_o;
    reg [63:0] l_TColl_0_2_2_constprop_o;
    reg [63:0] l_TColl_0_2_3_constprop_o;
    reg [63:0] l_TColl_1_2_0_constprop_o;
    reg [63:0] l_TColl_1_2_1_constprop_o;
    reg [63:0] l_TColl_1_2_2_constprop_o;
    reg [63:0] l_TColl_1_2_3_constprop_o;
    reg [63:0] l_TColl_2_2_0_constprop_o;
    reg [63:0] l_TColl_2_2_1_constprop_o;
    reg [63:0] l_TColl_2_2_2_constprop_o;
    reg [63:0] l_TColl_2_2_3_constprop_o;
    reg [63:0] l_TColl_0_3_0_constprop_o;
    reg [63:0] l_TColl_0_3_1_constprop_o;
    reg [63:0] l_TColl_0_3_2_constprop_o;
    reg [63:0] l_TColl_0_3_3_constprop_o;
    reg [63:0] l_TColl_1_3_0_constprop_o;
    reg [63:0] l_TColl_1_3_1_constprop_o;
    reg [63:0] l_TColl_1_3_2_constprop_o;
    reg [63:0] l_TColl_1_3_3_constprop_o;
    reg [63:0] l_TColl_2_3_0_constprop_o;
    reg [63:0] l_TColl_2_3_1_constprop_o;
    reg [63:0] l_TColl_2_3_2_constprop_o;
    reg [63:0] l_TColl_2_3_3_constprop_o;
    reg [0:0] ap_return;

    (* fsm_encoding = "none" *) reg [7:0] ap_CS_fsm;
    wire ap_CS_fsm_state1;
    wire ap_CS_fsm_state3;
    wire [2:0] add_ln168_fu_1333_p2;
    reg [2:0] add_ln168_reg_1721;
    wire ap_CS_fsm_state5;
    wire [1:0] trunc_ln168_fu_1339_p1;
    reg [1:0] trunc_ln168_reg_1726;
    wire [4:0] tmp_48_fu_1343_p3;
    reg [4:0] tmp_48_reg_1731;
    wire [3:0] add_ln169_fu_1357_p2;
    reg [3:0] add_ln169_reg_1739;
    wire ap_CS_fsm_state6;
    wire [2:0] trunc_ln169_fu_1367_p1;
    reg [2:0] trunc_ln169_reg_1744;
    wire [4:0] add_ln170_fu_1372_p2;
    reg [4:0] add_ln170_reg_1749;
    reg [4:0] checks_address0;
    reg checks_ce0;
    reg checks_we0;
    reg [0:0] checks_d0;
    wire [0:0] checks_q0;
    wire grp_forwardKin_fu_863_ap_start;
    wire grp_forwardKin_fu_863_ap_done;
    wire grp_forwardKin_fu_863_ap_idle;
    wire grp_forwardKin_fu_863_ap_ready;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_0_0_address0;
    wire grp_forwardKin_fu_863_this_TLink_0_0_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_0_1_address0;
    wire grp_forwardKin_fu_863_this_TLink_0_1_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_0_2_address0;
    wire grp_forwardKin_fu_863_this_TLink_0_2_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_0_3_address0;
    wire grp_forwardKin_fu_863_this_TLink_0_3_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_1_0_address0;
    wire grp_forwardKin_fu_863_this_TLink_1_0_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_1_1_address0;
    wire grp_forwardKin_fu_863_this_TLink_1_1_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_1_2_address0;
    wire grp_forwardKin_fu_863_this_TLink_1_2_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_1_3_address0;
    wire grp_forwardKin_fu_863_this_TLink_1_3_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_2_0_address0;
    wire grp_forwardKin_fu_863_this_TLink_2_0_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_2_1_address0;
    wire grp_forwardKin_fu_863_this_TLink_2_1_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_2_2_address0;
    wire grp_forwardKin_fu_863_this_TLink_2_2_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_2_3_address0;
    wire grp_forwardKin_fu_863_this_TLink_2_3_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_3_0_address0;
    wire grp_forwardKin_fu_863_this_TLink_3_0_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_3_1_address0;
    wire grp_forwardKin_fu_863_this_TLink_3_1_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_3_2_address0;
    wire grp_forwardKin_fu_863_this_TLink_3_2_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TLink_3_3_address0;
    wire grp_forwardKin_fu_863_this_TLink_3_3_ce0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_0_0_address0;
    wire grp_forwardKin_fu_863_this_TJoint_0_0_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_0_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_0_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_0_1_address0;
    wire grp_forwardKin_fu_863_this_TJoint_0_1_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_0_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_0_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_0_2_address0;
    wire grp_forwardKin_fu_863_this_TJoint_0_2_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_0_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_0_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_0_3_address0;
    wire grp_forwardKin_fu_863_this_TJoint_0_3_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_0_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_0_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_1_0_address0;
    wire grp_forwardKin_fu_863_this_TJoint_1_0_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_1_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_1_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_1_1_address0;
    wire grp_forwardKin_fu_863_this_TJoint_1_1_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_1_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_1_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_1_2_address0;
    wire grp_forwardKin_fu_863_this_TJoint_1_2_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_1_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_1_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_1_3_address0;
    wire grp_forwardKin_fu_863_this_TJoint_1_3_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_1_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_1_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_2_0_address0;
    wire grp_forwardKin_fu_863_this_TJoint_2_0_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_2_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_2_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_2_1_address0;
    wire grp_forwardKin_fu_863_this_TJoint_2_1_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_2_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_2_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_2_2_address0;
    wire grp_forwardKin_fu_863_this_TJoint_2_2_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_2_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_2_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_2_3_address0;
    wire grp_forwardKin_fu_863_this_TJoint_2_3_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_2_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_2_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_3_0_address0;
    wire grp_forwardKin_fu_863_this_TJoint_3_0_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_3_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_3_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_3_1_address0;
    wire grp_forwardKin_fu_863_this_TJoint_3_1_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_3_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_3_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_3_2_address0;
    wire grp_forwardKin_fu_863_this_TJoint_3_2_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_3_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_3_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TJoint_3_3_address0;
    wire grp_forwardKin_fu_863_this_TJoint_3_3_ce0;
    wire grp_forwardKin_fu_863_this_TJoint_3_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TJoint_3_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_0_0_address0;
    wire grp_forwardKin_fu_863_this_TCurr_0_0_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_0_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_0_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_0_1_address0;
    wire grp_forwardKin_fu_863_this_TCurr_0_1_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_0_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_0_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_0_2_address0;
    wire grp_forwardKin_fu_863_this_TCurr_0_2_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_0_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_0_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_0_3_address0;
    wire grp_forwardKin_fu_863_this_TCurr_0_3_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_0_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_0_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_1_0_address0;
    wire grp_forwardKin_fu_863_this_TCurr_1_0_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_1_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_1_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_1_1_address0;
    wire grp_forwardKin_fu_863_this_TCurr_1_1_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_1_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_1_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_1_2_address0;
    wire grp_forwardKin_fu_863_this_TCurr_1_2_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_1_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_1_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_1_3_address0;
    wire grp_forwardKin_fu_863_this_TCurr_1_3_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_1_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_1_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_2_0_address0;
    wire grp_forwardKin_fu_863_this_TCurr_2_0_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_2_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_2_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_2_1_address0;
    wire grp_forwardKin_fu_863_this_TCurr_2_1_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_2_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_2_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_2_2_address0;
    wire grp_forwardKin_fu_863_this_TCurr_2_2_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_2_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_2_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_2_3_address0;
    wire grp_forwardKin_fu_863_this_TCurr_2_3_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_2_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_2_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_3_0_address0;
    wire grp_forwardKin_fu_863_this_TCurr_3_0_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_3_0_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_3_0_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_3_1_address0;
    wire grp_forwardKin_fu_863_this_TCurr_3_1_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_3_1_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_3_1_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_3_2_address0;
    wire grp_forwardKin_fu_863_this_TCurr_3_2_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_3_2_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_3_2_d0;
    wire [2:0] grp_forwardKin_fu_863_this_TCurr_3_3_address0;
    wire grp_forwardKin_fu_863_this_TCurr_3_3_ce0;
    wire grp_forwardKin_fu_863_this_TCurr_3_3_we0;
    wire [63:0] grp_forwardKin_fu_863_this_TCurr_3_3_d0;
    wire [2:0] grp_forwardKin_fu_863_this_q_address0;
    wire grp_forwardKin_fu_863_this_q_ce0;
    wire grp_forwardKin_fu_863_this_q_we0;
    wire [63:0] grp_forwardKin_fu_863_this_q_d0;
    wire [2:0] grp_forwardKin_fu_863_ang_address0;
    wire grp_forwardKin_fu_863_ang_ce0;
    wire grp_detectCollNode_Pipeline_2_fu_985_ap_start;
    wire grp_detectCollNode_Pipeline_2_fu_985_ap_done;
    wire grp_detectCollNode_Pipeline_2_fu_985_ap_idle;
    wire grp_detectCollNode_Pipeline_2_fu_985_ap_ready;
    wire [4:0] grp_detectCollNode_Pipeline_2_fu_985_checks_address0;
    wire grp_detectCollNode_Pipeline_2_fu_985_checks_ce0;
    wire grp_detectCollNode_Pipeline_2_fu_985_checks_we0;
    wire [0:0] grp_detectCollNode_Pipeline_2_fu_985_checks_d0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_done;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_idle;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_ready;
    wire [6:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we0;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d0;
    wire [6:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address1;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce1;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we1;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d1;
    wire [5:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_ce0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_we0;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_d0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_ce0;
    wire [2:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_ce0;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din0;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din1;
    wire [0:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_opcode;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_ce;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din0;
    wire [63:0] grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din1;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_ce;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_idle;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_ready;
    wire [4:0] grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_address0;
    wire grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_ce0;
    wire [0:0] grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_return;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_ap_start;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_ap_done;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_ap_idle;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_ap_ready;
    wire [6:0] grp_cuboidCuboidCollision_double_s_fu_1252_p1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_s_fu_1252_p1_address1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce1;
    wire [5:0] grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce0;
    wire [5:0] grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce1;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_ce0;
    wire [2:0] grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address0;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce0;
    wire [6:0] grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce1;
    wire [0:0] grp_cuboidCuboidCollision_double_s_fu_1252_ap_return;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din1;
    wire [1:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din1;
    wire [4:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_opcode;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_ce;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din0;
    wire [63:0] grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din1;
    wire grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_ce;
    reg [3:0] j_reg_852;
    wire ap_CS_fsm_state7;
    wire [0:0] icmp_ln168_fu_1327_p2;
    reg grp_forwardKin_fu_863_ap_start_reg;
    wire ap_CS_fsm_state2;
    reg grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg;
    reg grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg;
    wire ap_CS_fsm_state4;
    reg grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg;
    wire ap_CS_fsm_state8;
    reg grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg;
    wire [0:0] icmp_ln169_fu_1351_p2;
    wire [63:0] zext_ln170_fu_1381_p1;
    reg [2:0] i_fu_448;
    wire [4:0] zext_ln169_fu_1363_p1;
    wire [0:0] xor_ln176_fu_1385_p2;
    reg [63:0] grp_fu_1754_p0;
    reg [63:0] grp_fu_1754_p1;
    reg [1:0] grp_fu_1754_opcode;
    reg grp_fu_1754_ce;
    reg [63:0] grp_fu_1758_p0;
    reg [63:0] grp_fu_1758_p1;
    reg grp_fu_1758_ce;
    reg grp_fu_1762_ce;
    reg grp_fu_1766_ce;
    reg grp_fu_1770_ce;
    reg grp_fu_1774_ce;
    reg grp_fu_1778_ce;
    reg grp_fu_1782_ce;
    reg grp_fu_1786_ce;
    reg grp_fu_1790_ce;
    reg grp_fu_1794_ce;
    reg grp_fu_1798_ce;
    reg [0:0] ap_return_preg;
    reg [7:0] ap_NS_fsm;
    reg ap_ST_fsm_state1_blk;
    reg ap_block_state2_on_subcall_done;
    reg ap_ST_fsm_state2_blk;
    wire ap_ST_fsm_state3_blk;
    reg ap_ST_fsm_state4_blk;
    wire ap_ST_fsm_state5_blk;
    wire ap_ST_fsm_state6_blk;
    reg ap_ST_fsm_state7_blk;
    reg ap_ST_fsm_state8_blk;
    wire ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 8'd1;
        #0 grp_forwardKin_fu_863_ap_start_reg = 1'b0;
        #0 grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg = 1'b0;
        #0 grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg = 1'b0;
        #0 grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg = 1'b0;
        #0 grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg = 1'b0;
        #0 i_fu_448 = 3'd0;
        #0 ap_return_preg = 1'd0;
    end

    main_detectCollNode_checks_RAM_AUTO_1R1W #(
        .DataWidth(1),
        .AddressRange(32),
        .AddressWidth(5)
    ) checks_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(checks_address0),
        .ce0(checks_ce0),
        .we0(checks_we0),
        .d0(checks_d0),
        .q0(checks_q0)
    );

    main_forwardKin grp_forwardKin_fu_863 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_forwardKin_fu_863_ap_start),
        .ap_done(grp_forwardKin_fu_863_ap_done),
        .ap_idle(grp_forwardKin_fu_863_ap_idle),
        .ap_ready(grp_forwardKin_fu_863_ap_ready),
        .this_TLink_0_0_address0(grp_forwardKin_fu_863_this_TLink_0_0_address0),
        .this_TLink_0_0_ce0(grp_forwardKin_fu_863_this_TLink_0_0_ce0),
        .this_TLink_0_0_q0(this_TLink_0_0_q0),
        .this_TLink_0_1_address0(grp_forwardKin_fu_863_this_TLink_0_1_address0),
        .this_TLink_0_1_ce0(grp_forwardKin_fu_863_this_TLink_0_1_ce0),
        .this_TLink_0_1_q0(this_TLink_0_1_q0),
        .this_TLink_0_2_address0(grp_forwardKin_fu_863_this_TLink_0_2_address0),
        .this_TLink_0_2_ce0(grp_forwardKin_fu_863_this_TLink_0_2_ce0),
        .this_TLink_0_2_q0(this_TLink_0_2_q0),
        .this_TLink_0_3_address0(grp_forwardKin_fu_863_this_TLink_0_3_address0),
        .this_TLink_0_3_ce0(grp_forwardKin_fu_863_this_TLink_0_3_ce0),
        .this_TLink_0_3_q0(this_TLink_0_3_q0),
        .this_TLink_1_0_address0(grp_forwardKin_fu_863_this_TLink_1_0_address0),
        .this_TLink_1_0_ce0(grp_forwardKin_fu_863_this_TLink_1_0_ce0),
        .this_TLink_1_0_q0(this_TLink_1_0_q0),
        .this_TLink_1_1_address0(grp_forwardKin_fu_863_this_TLink_1_1_address0),
        .this_TLink_1_1_ce0(grp_forwardKin_fu_863_this_TLink_1_1_ce0),
        .this_TLink_1_1_q0(this_TLink_1_1_q0),
        .this_TLink_1_2_address0(grp_forwardKin_fu_863_this_TLink_1_2_address0),
        .this_TLink_1_2_ce0(grp_forwardKin_fu_863_this_TLink_1_2_ce0),
        .this_TLink_1_2_q0(this_TLink_1_2_q0),
        .this_TLink_1_3_address0(grp_forwardKin_fu_863_this_TLink_1_3_address0),
        .this_TLink_1_3_ce0(grp_forwardKin_fu_863_this_TLink_1_3_ce0),
        .this_TLink_1_3_q0(this_TLink_1_3_q0),
        .this_TLink_2_0_address0(grp_forwardKin_fu_863_this_TLink_2_0_address0),
        .this_TLink_2_0_ce0(grp_forwardKin_fu_863_this_TLink_2_0_ce0),
        .this_TLink_2_0_q0(this_TLink_2_0_q0),
        .this_TLink_2_1_address0(grp_forwardKin_fu_863_this_TLink_2_1_address0),
        .this_TLink_2_1_ce0(grp_forwardKin_fu_863_this_TLink_2_1_ce0),
        .this_TLink_2_1_q0(this_TLink_2_1_q0),
        .this_TLink_2_2_address0(grp_forwardKin_fu_863_this_TLink_2_2_address0),
        .this_TLink_2_2_ce0(grp_forwardKin_fu_863_this_TLink_2_2_ce0),
        .this_TLink_2_2_q0(this_TLink_2_2_q0),
        .this_TLink_2_3_address0(grp_forwardKin_fu_863_this_TLink_2_3_address0),
        .this_TLink_2_3_ce0(grp_forwardKin_fu_863_this_TLink_2_3_ce0),
        .this_TLink_2_3_q0(this_TLink_2_3_q0),
        .this_TLink_3_0_address0(grp_forwardKin_fu_863_this_TLink_3_0_address0),
        .this_TLink_3_0_ce0(grp_forwardKin_fu_863_this_TLink_3_0_ce0),
        .this_TLink_3_0_q0(this_TLink_3_0_q0),
        .this_TLink_3_1_address0(grp_forwardKin_fu_863_this_TLink_3_1_address0),
        .this_TLink_3_1_ce0(grp_forwardKin_fu_863_this_TLink_3_1_ce0),
        .this_TLink_3_1_q0(this_TLink_3_1_q0),
        .this_TLink_3_2_address0(grp_forwardKin_fu_863_this_TLink_3_2_address0),
        .this_TLink_3_2_ce0(grp_forwardKin_fu_863_this_TLink_3_2_ce0),
        .this_TLink_3_2_q0(this_TLink_3_2_q0),
        .this_TLink_3_3_address0(grp_forwardKin_fu_863_this_TLink_3_3_address0),
        .this_TLink_3_3_ce0(grp_forwardKin_fu_863_this_TLink_3_3_ce0),
        .this_TLink_3_3_q0(this_TLink_3_3_q0),
        .this_TJoint_0_0_address0(grp_forwardKin_fu_863_this_TJoint_0_0_address0),
        .this_TJoint_0_0_ce0(grp_forwardKin_fu_863_this_TJoint_0_0_ce0),
        .this_TJoint_0_0_we0(grp_forwardKin_fu_863_this_TJoint_0_0_we0),
        .this_TJoint_0_0_d0(grp_forwardKin_fu_863_this_TJoint_0_0_d0),
        .this_TJoint_0_0_q0(this_TJoint_0_0_q0),
        .this_TJoint_0_1_address0(grp_forwardKin_fu_863_this_TJoint_0_1_address0),
        .this_TJoint_0_1_ce0(grp_forwardKin_fu_863_this_TJoint_0_1_ce0),
        .this_TJoint_0_1_we0(grp_forwardKin_fu_863_this_TJoint_0_1_we0),
        .this_TJoint_0_1_d0(grp_forwardKin_fu_863_this_TJoint_0_1_d0),
        .this_TJoint_0_1_q0(this_TJoint_0_1_q0),
        .this_TJoint_0_2_address0(grp_forwardKin_fu_863_this_TJoint_0_2_address0),
        .this_TJoint_0_2_ce0(grp_forwardKin_fu_863_this_TJoint_0_2_ce0),
        .this_TJoint_0_2_we0(grp_forwardKin_fu_863_this_TJoint_0_2_we0),
        .this_TJoint_0_2_d0(grp_forwardKin_fu_863_this_TJoint_0_2_d0),
        .this_TJoint_0_2_q0(this_TJoint_0_2_q0),
        .this_TJoint_0_3_address0(grp_forwardKin_fu_863_this_TJoint_0_3_address0),
        .this_TJoint_0_3_ce0(grp_forwardKin_fu_863_this_TJoint_0_3_ce0),
        .this_TJoint_0_3_we0(grp_forwardKin_fu_863_this_TJoint_0_3_we0),
        .this_TJoint_0_3_d0(grp_forwardKin_fu_863_this_TJoint_0_3_d0),
        .this_TJoint_0_3_q0(this_TJoint_0_3_q0),
        .this_TJoint_1_0_address0(grp_forwardKin_fu_863_this_TJoint_1_0_address0),
        .this_TJoint_1_0_ce0(grp_forwardKin_fu_863_this_TJoint_1_0_ce0),
        .this_TJoint_1_0_we0(grp_forwardKin_fu_863_this_TJoint_1_0_we0),
        .this_TJoint_1_0_d0(grp_forwardKin_fu_863_this_TJoint_1_0_d0),
        .this_TJoint_1_0_q0(this_TJoint_1_0_q0),
        .this_TJoint_1_1_address0(grp_forwardKin_fu_863_this_TJoint_1_1_address0),
        .this_TJoint_1_1_ce0(grp_forwardKin_fu_863_this_TJoint_1_1_ce0),
        .this_TJoint_1_1_we0(grp_forwardKin_fu_863_this_TJoint_1_1_we0),
        .this_TJoint_1_1_d0(grp_forwardKin_fu_863_this_TJoint_1_1_d0),
        .this_TJoint_1_1_q0(this_TJoint_1_1_q0),
        .this_TJoint_1_2_address0(grp_forwardKin_fu_863_this_TJoint_1_2_address0),
        .this_TJoint_1_2_ce0(grp_forwardKin_fu_863_this_TJoint_1_2_ce0),
        .this_TJoint_1_2_we0(grp_forwardKin_fu_863_this_TJoint_1_2_we0),
        .this_TJoint_1_2_d0(grp_forwardKin_fu_863_this_TJoint_1_2_d0),
        .this_TJoint_1_2_q0(this_TJoint_1_2_q0),
        .this_TJoint_1_3_address0(grp_forwardKin_fu_863_this_TJoint_1_3_address0),
        .this_TJoint_1_3_ce0(grp_forwardKin_fu_863_this_TJoint_1_3_ce0),
        .this_TJoint_1_3_we0(grp_forwardKin_fu_863_this_TJoint_1_3_we0),
        .this_TJoint_1_3_d0(grp_forwardKin_fu_863_this_TJoint_1_3_d0),
        .this_TJoint_1_3_q0(this_TJoint_1_3_q0),
        .this_TJoint_2_0_address0(grp_forwardKin_fu_863_this_TJoint_2_0_address0),
        .this_TJoint_2_0_ce0(grp_forwardKin_fu_863_this_TJoint_2_0_ce0),
        .this_TJoint_2_0_we0(grp_forwardKin_fu_863_this_TJoint_2_0_we0),
        .this_TJoint_2_0_d0(grp_forwardKin_fu_863_this_TJoint_2_0_d0),
        .this_TJoint_2_0_q0(this_TJoint_2_0_q0),
        .this_TJoint_2_1_address0(grp_forwardKin_fu_863_this_TJoint_2_1_address0),
        .this_TJoint_2_1_ce0(grp_forwardKin_fu_863_this_TJoint_2_1_ce0),
        .this_TJoint_2_1_we0(grp_forwardKin_fu_863_this_TJoint_2_1_we0),
        .this_TJoint_2_1_d0(grp_forwardKin_fu_863_this_TJoint_2_1_d0),
        .this_TJoint_2_1_q0(this_TJoint_2_1_q0),
        .this_TJoint_2_2_address0(grp_forwardKin_fu_863_this_TJoint_2_2_address0),
        .this_TJoint_2_2_ce0(grp_forwardKin_fu_863_this_TJoint_2_2_ce0),
        .this_TJoint_2_2_we0(grp_forwardKin_fu_863_this_TJoint_2_2_we0),
        .this_TJoint_2_2_d0(grp_forwardKin_fu_863_this_TJoint_2_2_d0),
        .this_TJoint_2_2_q0(this_TJoint_2_2_q0),
        .this_TJoint_2_3_address0(grp_forwardKin_fu_863_this_TJoint_2_3_address0),
        .this_TJoint_2_3_ce0(grp_forwardKin_fu_863_this_TJoint_2_3_ce0),
        .this_TJoint_2_3_we0(grp_forwardKin_fu_863_this_TJoint_2_3_we0),
        .this_TJoint_2_3_d0(grp_forwardKin_fu_863_this_TJoint_2_3_d0),
        .this_TJoint_2_3_q0(this_TJoint_2_3_q0),
        .this_TJoint_3_0_address0(grp_forwardKin_fu_863_this_TJoint_3_0_address0),
        .this_TJoint_3_0_ce0(grp_forwardKin_fu_863_this_TJoint_3_0_ce0),
        .this_TJoint_3_0_we0(grp_forwardKin_fu_863_this_TJoint_3_0_we0),
        .this_TJoint_3_0_d0(grp_forwardKin_fu_863_this_TJoint_3_0_d0),
        .this_TJoint_3_0_q0(this_TJoint_3_0_q0),
        .this_TJoint_3_1_address0(grp_forwardKin_fu_863_this_TJoint_3_1_address0),
        .this_TJoint_3_1_ce0(grp_forwardKin_fu_863_this_TJoint_3_1_ce0),
        .this_TJoint_3_1_we0(grp_forwardKin_fu_863_this_TJoint_3_1_we0),
        .this_TJoint_3_1_d0(grp_forwardKin_fu_863_this_TJoint_3_1_d0),
        .this_TJoint_3_1_q0(this_TJoint_3_1_q0),
        .this_TJoint_3_2_address0(grp_forwardKin_fu_863_this_TJoint_3_2_address0),
        .this_TJoint_3_2_ce0(grp_forwardKin_fu_863_this_TJoint_3_2_ce0),
        .this_TJoint_3_2_we0(grp_forwardKin_fu_863_this_TJoint_3_2_we0),
        .this_TJoint_3_2_d0(grp_forwardKin_fu_863_this_TJoint_3_2_d0),
        .this_TJoint_3_2_q0(this_TJoint_3_2_q0),
        .this_TJoint_3_3_address0(grp_forwardKin_fu_863_this_TJoint_3_3_address0),
        .this_TJoint_3_3_ce0(grp_forwardKin_fu_863_this_TJoint_3_3_ce0),
        .this_TJoint_3_3_we0(grp_forwardKin_fu_863_this_TJoint_3_3_we0),
        .this_TJoint_3_3_d0(grp_forwardKin_fu_863_this_TJoint_3_3_d0),
        .this_TJoint_3_3_q0(this_TJoint_3_3_q0),
        .this_TCurr_0_0_address0(grp_forwardKin_fu_863_this_TCurr_0_0_address0),
        .this_TCurr_0_0_ce0(grp_forwardKin_fu_863_this_TCurr_0_0_ce0),
        .this_TCurr_0_0_we0(grp_forwardKin_fu_863_this_TCurr_0_0_we0),
        .this_TCurr_0_0_d0(grp_forwardKin_fu_863_this_TCurr_0_0_d0),
        .this_TCurr_0_0_q0(this_TCurr_0_0_q0),
        .this_TCurr_0_1_address0(grp_forwardKin_fu_863_this_TCurr_0_1_address0),
        .this_TCurr_0_1_ce0(grp_forwardKin_fu_863_this_TCurr_0_1_ce0),
        .this_TCurr_0_1_we0(grp_forwardKin_fu_863_this_TCurr_0_1_we0),
        .this_TCurr_0_1_d0(grp_forwardKin_fu_863_this_TCurr_0_1_d0),
        .this_TCurr_0_1_q0(this_TCurr_0_1_q0),
        .this_TCurr_0_2_address0(grp_forwardKin_fu_863_this_TCurr_0_2_address0),
        .this_TCurr_0_2_ce0(grp_forwardKin_fu_863_this_TCurr_0_2_ce0),
        .this_TCurr_0_2_we0(grp_forwardKin_fu_863_this_TCurr_0_2_we0),
        .this_TCurr_0_2_d0(grp_forwardKin_fu_863_this_TCurr_0_2_d0),
        .this_TCurr_0_2_q0(this_TCurr_0_2_q0),
        .this_TCurr_0_3_address0(grp_forwardKin_fu_863_this_TCurr_0_3_address0),
        .this_TCurr_0_3_ce0(grp_forwardKin_fu_863_this_TCurr_0_3_ce0),
        .this_TCurr_0_3_we0(grp_forwardKin_fu_863_this_TCurr_0_3_we0),
        .this_TCurr_0_3_d0(grp_forwardKin_fu_863_this_TCurr_0_3_d0),
        .this_TCurr_0_3_q0(this_TCurr_0_3_q0),
        .this_TCurr_1_0_address0(grp_forwardKin_fu_863_this_TCurr_1_0_address0),
        .this_TCurr_1_0_ce0(grp_forwardKin_fu_863_this_TCurr_1_0_ce0),
        .this_TCurr_1_0_we0(grp_forwardKin_fu_863_this_TCurr_1_0_we0),
        .this_TCurr_1_0_d0(grp_forwardKin_fu_863_this_TCurr_1_0_d0),
        .this_TCurr_1_0_q0(this_TCurr_1_0_q0),
        .this_TCurr_1_1_address0(grp_forwardKin_fu_863_this_TCurr_1_1_address0),
        .this_TCurr_1_1_ce0(grp_forwardKin_fu_863_this_TCurr_1_1_ce0),
        .this_TCurr_1_1_we0(grp_forwardKin_fu_863_this_TCurr_1_1_we0),
        .this_TCurr_1_1_d0(grp_forwardKin_fu_863_this_TCurr_1_1_d0),
        .this_TCurr_1_1_q0(this_TCurr_1_1_q0),
        .this_TCurr_1_2_address0(grp_forwardKin_fu_863_this_TCurr_1_2_address0),
        .this_TCurr_1_2_ce0(grp_forwardKin_fu_863_this_TCurr_1_2_ce0),
        .this_TCurr_1_2_we0(grp_forwardKin_fu_863_this_TCurr_1_2_we0),
        .this_TCurr_1_2_d0(grp_forwardKin_fu_863_this_TCurr_1_2_d0),
        .this_TCurr_1_2_q0(this_TCurr_1_2_q0),
        .this_TCurr_1_3_address0(grp_forwardKin_fu_863_this_TCurr_1_3_address0),
        .this_TCurr_1_3_ce0(grp_forwardKin_fu_863_this_TCurr_1_3_ce0),
        .this_TCurr_1_3_we0(grp_forwardKin_fu_863_this_TCurr_1_3_we0),
        .this_TCurr_1_3_d0(grp_forwardKin_fu_863_this_TCurr_1_3_d0),
        .this_TCurr_1_3_q0(this_TCurr_1_3_q0),
        .this_TCurr_2_0_address0(grp_forwardKin_fu_863_this_TCurr_2_0_address0),
        .this_TCurr_2_0_ce0(grp_forwardKin_fu_863_this_TCurr_2_0_ce0),
        .this_TCurr_2_0_we0(grp_forwardKin_fu_863_this_TCurr_2_0_we0),
        .this_TCurr_2_0_d0(grp_forwardKin_fu_863_this_TCurr_2_0_d0),
        .this_TCurr_2_0_q0(this_TCurr_2_0_q0),
        .this_TCurr_2_1_address0(grp_forwardKin_fu_863_this_TCurr_2_1_address0),
        .this_TCurr_2_1_ce0(grp_forwardKin_fu_863_this_TCurr_2_1_ce0),
        .this_TCurr_2_1_we0(grp_forwardKin_fu_863_this_TCurr_2_1_we0),
        .this_TCurr_2_1_d0(grp_forwardKin_fu_863_this_TCurr_2_1_d0),
        .this_TCurr_2_1_q0(this_TCurr_2_1_q0),
        .this_TCurr_2_2_address0(grp_forwardKin_fu_863_this_TCurr_2_2_address0),
        .this_TCurr_2_2_ce0(grp_forwardKin_fu_863_this_TCurr_2_2_ce0),
        .this_TCurr_2_2_we0(grp_forwardKin_fu_863_this_TCurr_2_2_we0),
        .this_TCurr_2_2_d0(grp_forwardKin_fu_863_this_TCurr_2_2_d0),
        .this_TCurr_2_2_q0(this_TCurr_2_2_q0),
        .this_TCurr_2_3_address0(grp_forwardKin_fu_863_this_TCurr_2_3_address0),
        .this_TCurr_2_3_ce0(grp_forwardKin_fu_863_this_TCurr_2_3_ce0),
        .this_TCurr_2_3_we0(grp_forwardKin_fu_863_this_TCurr_2_3_we0),
        .this_TCurr_2_3_d0(grp_forwardKin_fu_863_this_TCurr_2_3_d0),
        .this_TCurr_2_3_q0(this_TCurr_2_3_q0),
        .this_TCurr_3_0_address0(grp_forwardKin_fu_863_this_TCurr_3_0_address0),
        .this_TCurr_3_0_ce0(grp_forwardKin_fu_863_this_TCurr_3_0_ce0),
        .this_TCurr_3_0_we0(grp_forwardKin_fu_863_this_TCurr_3_0_we0),
        .this_TCurr_3_0_d0(grp_forwardKin_fu_863_this_TCurr_3_0_d0),
        .this_TCurr_3_0_q0(this_TCurr_3_0_q0),
        .this_TCurr_3_1_address0(grp_forwardKin_fu_863_this_TCurr_3_1_address0),
        .this_TCurr_3_1_ce0(grp_forwardKin_fu_863_this_TCurr_3_1_ce0),
        .this_TCurr_3_1_we0(grp_forwardKin_fu_863_this_TCurr_3_1_we0),
        .this_TCurr_3_1_d0(grp_forwardKin_fu_863_this_TCurr_3_1_d0),
        .this_TCurr_3_1_q0(this_TCurr_3_1_q0),
        .this_TCurr_3_2_address0(grp_forwardKin_fu_863_this_TCurr_3_2_address0),
        .this_TCurr_3_2_ce0(grp_forwardKin_fu_863_this_TCurr_3_2_ce0),
        .this_TCurr_3_2_we0(grp_forwardKin_fu_863_this_TCurr_3_2_we0),
        .this_TCurr_3_2_d0(grp_forwardKin_fu_863_this_TCurr_3_2_d0),
        .this_TCurr_3_2_q0(this_TCurr_3_2_q0),
        .this_TCurr_3_3_address0(grp_forwardKin_fu_863_this_TCurr_3_3_address0),
        .this_TCurr_3_3_ce0(grp_forwardKin_fu_863_this_TCurr_3_3_ce0),
        .this_TCurr_3_3_we0(grp_forwardKin_fu_863_this_TCurr_3_3_we0),
        .this_TCurr_3_3_d0(grp_forwardKin_fu_863_this_TCurr_3_3_d0),
        .this_TCurr_3_3_q0(this_TCurr_3_3_q0),
        .this_q_address0(grp_forwardKin_fu_863_this_q_address0),
        .this_q_ce0(grp_forwardKin_fu_863_this_q_ce0),
        .this_q_we0(grp_forwardKin_fu_863_this_q_we0),
        .this_q_d0(grp_forwardKin_fu_863_this_q_d0),
        .this_q_q0(this_q_q0),
        .ang_address0(grp_forwardKin_fu_863_ang_address0),
        .ang_ce0(grp_forwardKin_fu_863_ang_ce0),
        .ang_q0(ang_q0)
    );

    main_detectCollNode_Pipeline_2 grp_detectCollNode_Pipeline_2_fu_985 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_detectCollNode_Pipeline_2_fu_985_ap_start),
        .ap_done(grp_detectCollNode_Pipeline_2_fu_985_ap_done),
        .ap_idle(grp_detectCollNode_Pipeline_2_fu_985_ap_idle),
        .ap_ready(grp_detectCollNode_Pipeline_2_fu_985_ap_ready),
        .checks_address0(grp_detectCollNode_Pipeline_2_fu_985_checks_address0),
        .checks_ce0(grp_detectCollNode_Pipeline_2_fu_985_checks_ce0),
        .checks_we0(grp_detectCollNode_Pipeline_2_fu_985_checks_we0),
        .checks_d0(grp_detectCollNode_Pipeline_2_fu_985_checks_d0)
    );

    main_detectCollNode_Pipeline_VITIS_LOOP_276_1 grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start),
        .ap_done(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_done),
        .ap_idle(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_idle),
        .ap_ready(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_ready),
        .this_cPoints_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address0),
        .this_cPoints_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce0),
        .this_cPoints_we0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we0),
        .this_cPoints_d0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d0),
        .this_cPoints_address1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address1),
        .this_cPoints_ce1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce1),
        .this_cPoints_we1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we1),
        .this_cPoints_d1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d1),
        .this_cAxes_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_address0),
        .this_cAxes_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_ce0),
        .this_cAxes_we0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_we0),
        .this_cAxes_d0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_d0),
        .this_TCurr_0_0_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_address0),
        .this_TCurr_0_0_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_ce0),
        .this_TCurr_0_0_q0(this_TCurr_0_0_q0),
        .p_read(p_read),
        .p_read1(p_read1),
        .p_read2(p_read2),
        .p_read3(p_read3),
        .this_TCurr_0_1_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_address0),
        .this_TCurr_0_1_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_ce0),
        .this_TCurr_0_1_q0(this_TCurr_0_1_q0),
        .p_read16(p_read16),
        .p_read17(p_read17),
        .p_read18(p_read18),
        .p_read19(p_read19),
        .this_TCurr_0_2_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_address0),
        .this_TCurr_0_2_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_ce0),
        .this_TCurr_0_2_q0(this_TCurr_0_2_q0),
        .p_read32(p_read32),
        .p_read33(p_read33),
        .p_read34(p_read34),
        .p_read35(p_read35),
        .this_TCurr_0_3_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_address0),
        .this_TCurr_0_3_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_ce0),
        .this_TCurr_0_3_q0(this_TCurr_0_3_q0),
        .p_read48(p_read48),
        .p_read49(p_read49),
        .p_read50(p_read50),
        .p_read51(p_read51),
        .p_read4(p_read4),
        .p_read5(p_read5),
        .p_read6(p_read6),
        .p_read7(p_read7),
        .p_read20(p_read20),
        .p_read21(p_read21),
        .p_read22(p_read22),
        .p_read23(p_read23),
        .p_read36(p_read36),
        .p_read37(p_read37),
        .p_read38(p_read38),
        .p_read39(p_read39),
        .p_read52(p_read52),
        .p_read53(p_read53),
        .p_read54(p_read54),
        .p_read55(p_read55),
        .p_read8(p_read8),
        .p_read9(p_read9),
        .p_read10(p_read10),
        .p_read11(p_read11),
        .p_read24(p_read24),
        .p_read25(p_read25),
        .p_read26(p_read26),
        .p_read27(p_read27),
        .p_read40(p_read40),
        .p_read41(p_read41),
        .p_read42(p_read42),
        .p_read43(p_read43),
        .p_read56(p_read56),
        .p_read57(p_read57),
        .p_read58(p_read58),
        .p_read59(p_read59),
        .p_read12(p_read12),
        .p_read13(p_read13),
        .p_read14(p_read14),
        .p_read15(p_read15),
        .p_read28(p_read28),
        .p_read29(p_read29),
        .p_read30(p_read30),
        .p_read31(p_read31),
        .p_read44(p_read44),
        .p_read45(p_read45),
        .p_read46(p_read46),
        .p_read47(p_read47),
        .p_read60(p_read60),
        .p_read61(p_read61),
        .p_read62(p_read62),
        .p_read63(p_read63),
        .this_TCurr_1_0_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_address0),
        .this_TCurr_1_0_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_ce0),
        .this_TCurr_1_0_q0(this_TCurr_1_0_q0),
        .this_TCurr_1_1_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_address0),
        .this_TCurr_1_1_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_ce0),
        .this_TCurr_1_1_q0(this_TCurr_1_1_q0),
        .this_TCurr_1_2_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_address0),
        .this_TCurr_1_2_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_ce0),
        .this_TCurr_1_2_q0(this_TCurr_1_2_q0),
        .this_TCurr_1_3_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_address0),
        .this_TCurr_1_3_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_ce0),
        .this_TCurr_1_3_q0(this_TCurr_1_3_q0),
        .this_TCurr_2_0_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_address0),
        .this_TCurr_2_0_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_ce0),
        .this_TCurr_2_0_q0(this_TCurr_2_0_q0),
        .this_TCurr_2_1_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_address0),
        .this_TCurr_2_1_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_ce0),
        .this_TCurr_2_1_q0(this_TCurr_2_1_q0),
        .this_TCurr_2_2_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_address0),
        .this_TCurr_2_2_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_ce0),
        .this_TCurr_2_2_q0(this_TCurr_2_2_q0),
        .this_TCurr_2_3_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_address0),
        .this_TCurr_2_3_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_ce0),
        .this_TCurr_2_3_q0(this_TCurr_2_3_q0),
        .l_TColl_0_0_0_constprop_i(l_TColl_0_0_0_constprop_i),
        .l_TColl_0_0_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o),
        .l_TColl_0_0_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o_ap_vld),
        .l_TColl_0_0_1_constprop_i(l_TColl_0_0_1_constprop_i),
        .l_TColl_0_0_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o),
        .l_TColl_0_0_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o_ap_vld),
        .l_TColl_0_0_2_constprop_i(l_TColl_0_0_2_constprop_i),
        .l_TColl_0_0_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o),
        .l_TColl_0_0_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o_ap_vld),
        .l_TColl_0_0_3_constprop_i(l_TColl_0_0_3_constprop_i),
        .l_TColl_0_0_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o),
        .l_TColl_0_0_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o_ap_vld),
        .l_TColl_1_0_0_constprop_i(l_TColl_1_0_0_constprop_i),
        .l_TColl_1_0_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o),
        .l_TColl_1_0_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o_ap_vld),
        .l_TColl_1_0_1_constprop_i(l_TColl_1_0_1_constprop_i),
        .l_TColl_1_0_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o),
        .l_TColl_1_0_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o_ap_vld),
        .l_TColl_1_0_2_constprop_i(l_TColl_1_0_2_constprop_i),
        .l_TColl_1_0_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o),
        .l_TColl_1_0_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o_ap_vld),
        .l_TColl_1_0_3_constprop_i(l_TColl_1_0_3_constprop_i),
        .l_TColl_1_0_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o),
        .l_TColl_1_0_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o_ap_vld),
        .l_TColl_2_0_0_constprop_i(l_TColl_2_0_0_constprop_i),
        .l_TColl_2_0_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o),
        .l_TColl_2_0_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o_ap_vld),
        .l_TColl_2_0_1_constprop_i(l_TColl_2_0_1_constprop_i),
        .l_TColl_2_0_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o),
        .l_TColl_2_0_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o_ap_vld),
        .l_TColl_2_0_2_constprop_i(l_TColl_2_0_2_constprop_i),
        .l_TColl_2_0_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o),
        .l_TColl_2_0_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o_ap_vld),
        .l_TColl_2_0_3_constprop_i(l_TColl_2_0_3_constprop_i),
        .l_TColl_2_0_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o),
        .l_TColl_2_0_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o_ap_vld),
        .l_TColl_0_1_0_constprop_i(l_TColl_0_1_0_constprop_i),
        .l_TColl_0_1_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o),
        .l_TColl_0_1_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o_ap_vld),
        .l_TColl_0_1_1_constprop_i(l_TColl_0_1_1_constprop_i),
        .l_TColl_0_1_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o),
        .l_TColl_0_1_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o_ap_vld),
        .l_TColl_0_1_2_constprop_i(l_TColl_0_1_2_constprop_i),
        .l_TColl_0_1_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o),
        .l_TColl_0_1_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o_ap_vld),
        .l_TColl_0_1_3_constprop_i(l_TColl_0_1_3_constprop_i),
        .l_TColl_0_1_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o),
        .l_TColl_0_1_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o_ap_vld),
        .l_TColl_1_1_0_constprop_i(l_TColl_1_1_0_constprop_i),
        .l_TColl_1_1_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o),
        .l_TColl_1_1_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o_ap_vld),
        .l_TColl_1_1_1_constprop_i(l_TColl_1_1_1_constprop_i),
        .l_TColl_1_1_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o),
        .l_TColl_1_1_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o_ap_vld),
        .l_TColl_1_1_2_constprop_i(l_TColl_1_1_2_constprop_i),
        .l_TColl_1_1_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o),
        .l_TColl_1_1_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o_ap_vld),
        .l_TColl_1_1_3_constprop_i(l_TColl_1_1_3_constprop_i),
        .l_TColl_1_1_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o),
        .l_TColl_1_1_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o_ap_vld),
        .l_TColl_2_1_0_constprop_i(l_TColl_2_1_0_constprop_i),
        .l_TColl_2_1_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o),
        .l_TColl_2_1_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o_ap_vld),
        .l_TColl_2_1_1_constprop_i(l_TColl_2_1_1_constprop_i),
        .l_TColl_2_1_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o),
        .l_TColl_2_1_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o_ap_vld),
        .l_TColl_2_1_2_constprop_i(l_TColl_2_1_2_constprop_i),
        .l_TColl_2_1_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o),
        .l_TColl_2_1_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o_ap_vld),
        .l_TColl_2_1_3_constprop_i(l_TColl_2_1_3_constprop_i),
        .l_TColl_2_1_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o),
        .l_TColl_2_1_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o_ap_vld),
        .l_TColl_0_2_0_constprop_i(l_TColl_0_2_0_constprop_i),
        .l_TColl_0_2_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o),
        .l_TColl_0_2_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o_ap_vld),
        .l_TColl_0_2_1_constprop_i(l_TColl_0_2_1_constprop_i),
        .l_TColl_0_2_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o),
        .l_TColl_0_2_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o_ap_vld),
        .l_TColl_0_2_2_constprop_i(l_TColl_0_2_2_constprop_i),
        .l_TColl_0_2_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o),
        .l_TColl_0_2_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o_ap_vld),
        .l_TColl_0_2_3_constprop_i(l_TColl_0_2_3_constprop_i),
        .l_TColl_0_2_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o),
        .l_TColl_0_2_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o_ap_vld),
        .l_TColl_1_2_0_constprop_i(l_TColl_1_2_0_constprop_i),
        .l_TColl_1_2_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o),
        .l_TColl_1_2_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o_ap_vld),
        .l_TColl_1_2_1_constprop_i(l_TColl_1_2_1_constprop_i),
        .l_TColl_1_2_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o),
        .l_TColl_1_2_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o_ap_vld),
        .l_TColl_1_2_2_constprop_i(l_TColl_1_2_2_constprop_i),
        .l_TColl_1_2_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o),
        .l_TColl_1_2_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o_ap_vld),
        .l_TColl_1_2_3_constprop_i(l_TColl_1_2_3_constprop_i),
        .l_TColl_1_2_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o),
        .l_TColl_1_2_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o_ap_vld),
        .l_TColl_2_2_0_constprop_i(l_TColl_2_2_0_constprop_i),
        .l_TColl_2_2_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o),
        .l_TColl_2_2_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o_ap_vld),
        .l_TColl_2_2_1_constprop_i(l_TColl_2_2_1_constprop_i),
        .l_TColl_2_2_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o),
        .l_TColl_2_2_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o_ap_vld),
        .l_TColl_2_2_2_constprop_i(l_TColl_2_2_2_constprop_i),
        .l_TColl_2_2_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o),
        .l_TColl_2_2_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o_ap_vld),
        .l_TColl_2_2_3_constprop_i(l_TColl_2_2_3_constprop_i),
        .l_TColl_2_2_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o),
        .l_TColl_2_2_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o_ap_vld),
        .l_TColl_0_3_0_constprop_i(l_TColl_0_3_0_constprop_i),
        .l_TColl_0_3_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o),
        .l_TColl_0_3_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o_ap_vld),
        .l_TColl_0_3_1_constprop_i(l_TColl_0_3_1_constprop_i),
        .l_TColl_0_3_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o),
        .l_TColl_0_3_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o_ap_vld),
        .l_TColl_0_3_2_constprop_i(l_TColl_0_3_2_constprop_i),
        .l_TColl_0_3_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o),
        .l_TColl_0_3_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o_ap_vld),
        .l_TColl_0_3_3_constprop_i(l_TColl_0_3_3_constprop_i),
        .l_TColl_0_3_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o),
        .l_TColl_0_3_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o_ap_vld),
        .l_TColl_1_3_0_constprop_i(l_TColl_1_3_0_constprop_i),
        .l_TColl_1_3_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o),
        .l_TColl_1_3_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o_ap_vld),
        .l_TColl_1_3_1_constprop_i(l_TColl_1_3_1_constprop_i),
        .l_TColl_1_3_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o),
        .l_TColl_1_3_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o_ap_vld),
        .l_TColl_1_3_2_constprop_i(l_TColl_1_3_2_constprop_i),
        .l_TColl_1_3_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o),
        .l_TColl_1_3_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o_ap_vld),
        .l_TColl_1_3_3_constprop_i(l_TColl_1_3_3_constprop_i),
        .l_TColl_1_3_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o),
        .l_TColl_1_3_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o_ap_vld),
        .l_TColl_2_3_0_constprop_i(l_TColl_2_3_0_constprop_i),
        .l_TColl_2_3_0_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o),
        .l_TColl_2_3_0_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o_ap_vld),
        .l_TColl_2_3_1_constprop_i(l_TColl_2_3_1_constprop_i),
        .l_TColl_2_3_1_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o),
        .l_TColl_2_3_1_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o_ap_vld),
        .l_TColl_2_3_2_constprop_i(l_TColl_2_3_2_constprop_i),
        .l_TColl_2_3_2_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o),
        .l_TColl_2_3_2_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o_ap_vld),
        .l_TColl_2_3_3_constprop_i(l_TColl_2_3_3_constprop_i),
        .l_TColl_2_3_3_constprop_o(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o),
        .l_TColl_2_3_3_constprop_o_ap_vld(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o_ap_vld),
        .grp_fu_1754_p_din0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din0),
        .grp_fu_1754_p_din1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din1),
        .grp_fu_1754_p_opcode(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_opcode),
        .grp_fu_1754_p_dout0(grp_fu_2529_p_dout0),
        .grp_fu_1754_p_ce(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_ce),
        .grp_fu_1758_p_din0(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din0),
        .grp_fu_1758_p_din1(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din1),
        .grp_fu_1758_p_dout0(grp_fu_2533_p_dout0),
        .grp_fu_1758_p_ce(grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_ce)
    );

    main_detectCollNode_Pipeline_VITIS_LOOP_176_3 grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start),
        .ap_done(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done),
        .ap_idle(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_idle),
        .ap_ready(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_ready),
        .checks_q0(checks_q0),
        .checks_address0(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_address0),
        .checks_ce0(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_ce0),
        .ap_return(grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_return)
    );

    main_cuboidCuboidCollision_double_s grp_cuboidCuboidCollision_double_s_fu_1252 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_cuboidCuboidCollision_double_s_fu_1252_ap_start),
        .ap_done(grp_cuboidCuboidCollision_double_s_fu_1252_ap_done),
        .ap_idle(grp_cuboidCuboidCollision_double_s_fu_1252_ap_idle),
        .ap_ready(grp_cuboidCuboidCollision_double_s_fu_1252_ap_ready),
        .p1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p1_address0),
        .p1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce0),
        .p1_q0(this_cPoints_q0),
        .p1_address1(grp_cuboidCuboidCollision_double_s_fu_1252_p1_address1),
        .p1_ce1(grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce1),
        .p1_q1(this_cPoints_q1),
        .p1_offset(trunc_ln168_reg_1726),
        .axes1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address0),
        .axes1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce0),
        .axes1_q0(this_cAxes_q0),
        .axes1_address1(grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address1),
        .axes1_ce1(grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce1),
        .axes1_q1(this_cAxes_q1),
        .p2_0_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_address0),
        .p2_0_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_ce0),
        .p2_0_0_q0(this_env_0_0_0_q0),
        .p2_0_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_address0),
        .p2_0_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_ce0),
        .p2_0_1_q0(this_env_0_0_1_q0),
        .p2_0_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_address0),
        .p2_0_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_ce0),
        .p2_0_2_q0(this_env_0_0_2_q0),
        .p2_1_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_address0),
        .p2_1_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_ce0),
        .p2_1_0_q0(this_env_0_1_0_q0),
        .p2_1_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_address0),
        .p2_1_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_ce0),
        .p2_1_1_q0(this_env_0_1_1_q0),
        .p2_1_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_address0),
        .p2_1_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_ce0),
        .p2_1_2_q0(this_env_0_1_2_q0),
        .p2_2_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_address0),
        .p2_2_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_ce0),
        .p2_2_0_q0(this_env_0_2_0_q0),
        .p2_2_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_address0),
        .p2_2_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_ce0),
        .p2_2_1_q0(this_env_0_2_1_q0),
        .p2_2_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_address0),
        .p2_2_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_ce0),
        .p2_2_2_q0(this_env_0_2_2_q0),
        .p2_3_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_address0),
        .p2_3_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_ce0),
        .p2_3_0_q0(this_env_0_3_0_q0),
        .p2_3_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_address0),
        .p2_3_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_ce0),
        .p2_3_1_q0(this_env_0_3_1_q0),
        .p2_3_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_address0),
        .p2_3_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_ce0),
        .p2_3_2_q0(this_env_0_3_2_q0),
        .p2_4_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_address0),
        .p2_4_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_ce0),
        .p2_4_0_q0(this_env_0_4_0_q0),
        .p2_4_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_address0),
        .p2_4_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_ce0),
        .p2_4_1_q0(this_env_0_4_1_q0),
        .p2_4_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_address0),
        .p2_4_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_ce0),
        .p2_4_2_q0(this_env_0_4_2_q0),
        .p2_5_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_address0),
        .p2_5_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_ce0),
        .p2_5_0_q0(this_env_0_5_0_q0),
        .p2_5_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_address0),
        .p2_5_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_ce0),
        .p2_5_1_q0(this_env_0_5_1_q0),
        .p2_5_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_address0),
        .p2_5_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_ce0),
        .p2_5_2_q0(this_env_0_5_2_q0),
        .p2_6_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_address0),
        .p2_6_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_ce0),
        .p2_6_0_q0(this_env_0_6_0_q0),
        .p2_6_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_address0),
        .p2_6_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_ce0),
        .p2_6_1_q0(this_env_0_6_1_q0),
        .p2_6_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_address0),
        .p2_6_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_ce0),
        .p2_6_2_q0(this_env_0_6_2_q0),
        .p2_7_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_address0),
        .p2_7_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_ce0),
        .p2_7_0_q0(this_env_0_7_0_q0),
        .p2_7_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_address0),
        .p2_7_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_ce0),
        .p2_7_1_q0(this_env_0_7_1_q0),
        .p2_7_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_address0),
        .p2_7_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_ce0),
        .p2_7_2_q0(this_env_0_7_2_q0),
        .p2_8_0_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_address0),
        .p2_8_0_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_ce0),
        .p2_8_0_q0(this_env_0_8_0_q0),
        .p2_8_1_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_address0),
        .p2_8_1_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_ce0),
        .p2_8_1_q0(this_env_0_8_1_q0),
        .p2_8_2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_address0),
        .p2_8_2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_ce0),
        .p2_8_2_q0(this_env_0_8_2_q0),
        .p2_offset(trunc_ln169_reg_1744),
        .axes2_address0(grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address0),
        .axes2_ce0(grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce0),
        .axes2_q0(this_env_1_q0),
        .axes2_address1(grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address1),
        .axes2_ce1(grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce1),
        .axes2_q1(this_env_1_q1),
        .ap_return(grp_cuboidCuboidCollision_double_s_fu_1252_ap_return),
        .grp_fu_1754_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din0),
        .grp_fu_1754_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din1),
        .grp_fu_1754_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_opcode),
        .grp_fu_1754_p_dout0(grp_fu_2529_p_dout0),
        .grp_fu_1754_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_ce),
        .grp_fu_1762_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din0),
        .grp_fu_1762_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din1),
        .grp_fu_1762_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_opcode),
        .grp_fu_1762_p_dout0(grp_fu_2537_p_dout0),
        .grp_fu_1762_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_ce),
        .grp_fu_1766_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din0),
        .grp_fu_1766_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din1),
        .grp_fu_1766_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_opcode),
        .grp_fu_1766_p_dout0(grp_fu_2541_p_dout0),
        .grp_fu_1766_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_ce),
        .grp_fu_1770_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din0),
        .grp_fu_1770_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din1),
        .grp_fu_1770_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_opcode),
        .grp_fu_1770_p_dout0(grp_fu_2545_p_dout0),
        .grp_fu_1770_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_ce),
        .grp_fu_1774_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din0),
        .grp_fu_1774_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din1),
        .grp_fu_1774_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_opcode),
        .grp_fu_1774_p_dout0(grp_fu_2549_p_dout0),
        .grp_fu_1774_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_ce),
        .grp_fu_1778_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din0),
        .grp_fu_1778_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din1),
        .grp_fu_1778_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_opcode),
        .grp_fu_1778_p_dout0(grp_fu_2553_p_dout0),
        .grp_fu_1778_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_ce),
        .grp_fu_1758_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din0),
        .grp_fu_1758_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din1),
        .grp_fu_1758_p_dout0(grp_fu_2533_p_dout0),
        .grp_fu_1758_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_ce),
        .grp_fu_1782_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din0),
        .grp_fu_1782_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din1),
        .grp_fu_1782_p_dout0(grp_fu_2557_p_dout0),
        .grp_fu_1782_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_ce),
        .grp_fu_1786_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din0),
        .grp_fu_1786_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din1),
        .grp_fu_1786_p_dout0(grp_fu_2561_p_dout0),
        .grp_fu_1786_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_ce),
        .grp_fu_1790_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din0),
        .grp_fu_1790_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din1),
        .grp_fu_1790_p_dout0(grp_fu_2565_p_dout0),
        .grp_fu_1790_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_ce),
        .grp_fu_1794_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din0),
        .grp_fu_1794_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din1),
        .grp_fu_1794_p_opcode(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_opcode),
        .grp_fu_1794_p_dout0(grp_fu_1454_p_dout0),
        .grp_fu_1794_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_ce),
        .grp_fu_1798_p_din0(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din0),
        .grp_fu_1798_p_din1(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din1),
        .grp_fu_1798_p_dout0(grp_fu_1462_p_dout0),
        .grp_fu_1798_p_ce(grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_ce)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg <= 1'd0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state8) & (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b1))) begin
                ap_return_preg <= xor_ln176_fu_1385_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state6) & (icmp_ln169_fu_1351_p2 == 1'd0))) begin
                grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg <= 1'b1;
            end else if ((grp_cuboidCuboidCollision_double_s_fu_1252_ap_ready == 1'b1)) begin
                grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg <= 1'b1;
            end else if ((grp_detectCollNode_Pipeline_2_fu_985_ap_ready == 1'b1)) begin
                grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state5) & (icmp_ln168_fu_1327_p2 == 1'd1))) begin
                grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg <= 1'b1;
            end else if ((grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_ready == 1'b1)) begin
                grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg <= 1'b1;
            end else if ((grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_ready == 1'b1)) begin
                grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_forwardKin_fu_863_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                grp_forwardKin_fu_863_ap_start_reg <= 1'b1;
            end else if ((grp_forwardKin_fu_863_ap_ready == 1'b1)) begin
                grp_forwardKin_fu_863_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
            i_fu_448 <= 3'd0;
        end else if (((1'b1 == ap_CS_fsm_state6) & (icmp_ln169_fu_1351_p2 == 1'd1))) begin
            i_fu_448 <= add_ln168_reg_1721;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state5) & (icmp_ln168_fu_1327_p2 == 1'd0))) begin
            j_reg_852 <= 4'd0;
        end else if (((1'b1 == ap_CS_fsm_state7) & (grp_cuboidCuboidCollision_double_s_fu_1252_ap_done == 1'b1))) begin
            j_reg_852 <= add_ln169_reg_1739;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            add_ln168_reg_1721 <= add_ln168_fu_1333_p2;
            tmp_48_reg_1731[4 : 3] <= tmp_48_fu_1343_p3[4 : 3];
            trunc_ln168_reg_1726 <= trunc_ln168_fu_1339_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state6)) begin
            add_ln169_reg_1739   <= add_ln169_fu_1357_p2;
            add_ln170_reg_1749   <= add_ln170_fu_1372_p2;
            trunc_ln169_reg_1744 <= trunc_ln169_fu_1367_p1;
        end
    end

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_block_state2_on_subcall_done)) begin
            ap_ST_fsm_state2_blk = 1'b1;
        end else begin
            ap_ST_fsm_state2_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state3_blk = 1'b0;

    always @(*) begin
        if ((grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_done == 1'b0)) begin
            ap_ST_fsm_state4_blk = 1'b1;
        end else begin
            ap_ST_fsm_state4_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state5_blk = 1'b0;

    assign ap_ST_fsm_state6_blk = 1'b0;

    always @(*) begin
        if ((grp_cuboidCuboidCollision_double_s_fu_1252_ap_done == 1'b0)) begin
            ap_ST_fsm_state7_blk = 1'b1;
        end else begin
            ap_ST_fsm_state7_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b0)) begin
            ap_ST_fsm_state8_blk = 1'b1;
        end else begin
            ap_ST_fsm_state8_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)) | ((1'b1 == ap_CS_fsm_state8) & (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b1))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b1))) begin
            ap_return = xor_ln176_fu_1385_p2;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            checks_address0 = zext_ln170_fu_1381_p1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            checks_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            checks_address0 = grp_detectCollNode_Pipeline_2_fu_985_checks_address0;
        end else begin
            checks_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state7) & (grp_cuboidCuboidCollision_double_s_fu_1252_ap_done == 1'b1))) begin
            checks_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            checks_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_checks_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            checks_ce0 = grp_detectCollNode_Pipeline_2_fu_985_checks_ce0;
        end else begin
            checks_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            checks_d0 = grp_cuboidCuboidCollision_double_s_fu_1252_ap_return;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            checks_d0 = grp_detectCollNode_Pipeline_2_fu_985_checks_d0;
        end else begin
            checks_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state7) & (grp_cuboidCuboidCollision_double_s_fu_1252_ap_done == 1'b1))) begin
            checks_we0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            checks_we0 = grp_detectCollNode_Pipeline_2_fu_985_checks_we0;
        end else begin
            checks_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1754_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1754_ce = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_ce;
        end else begin
            grp_fu_1754_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1754_opcode = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1754_opcode = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_opcode;
        end else begin
            grp_fu_1754_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1754_p0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1754_p0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din0;
        end else begin
            grp_fu_1754_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1754_p1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1754_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1754_p1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1754_p_din1;
        end else begin
            grp_fu_1754_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1758_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1758_ce = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_ce;
        end else begin
            grp_fu_1758_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1758_p0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1758_p0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din0;
        end else begin
            grp_fu_1758_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1758_p1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1758_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1758_p1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_grp_fu_1758_p_din1;
        end else begin
            grp_fu_1758_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1762_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_ce;
        end else begin
            grp_fu_1762_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1766_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_ce;
        end else begin
            grp_fu_1766_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1770_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_ce;
        end else begin
            grp_fu_1770_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1774_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_ce;
        end else begin
            grp_fu_1774_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1778_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_ce;
        end else begin
            grp_fu_1778_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1782_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_ce;
        end else begin
            grp_fu_1782_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1786_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_ce;
        end else begin
            grp_fu_1786_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1790_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_ce;
        end else begin
            grp_fu_1790_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1794_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_ce;
        end else begin
            grp_fu_1794_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            grp_fu_1798_ce = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_ce;
        end else begin
            grp_fu_1798_ce = 1'b1;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_0_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o;
        end else begin
            l_TColl_0_0_0_constprop_o = l_TColl_0_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_0_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o;
        end else begin
            l_TColl_0_0_1_constprop_o = l_TColl_0_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_0_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o;
        end else begin
            l_TColl_0_0_2_constprop_o = l_TColl_0_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_0_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o;
        end else begin
            l_TColl_0_0_3_constprop_o = l_TColl_0_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_1_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o;
        end else begin
            l_TColl_0_1_0_constprop_o = l_TColl_0_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_1_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o;
        end else begin
            l_TColl_0_1_1_constprop_o = l_TColl_0_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_1_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o;
        end else begin
            l_TColl_0_1_2_constprop_o = l_TColl_0_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_1_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o;
        end else begin
            l_TColl_0_1_3_constprop_o = l_TColl_0_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_2_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o;
        end else begin
            l_TColl_0_2_0_constprop_o = l_TColl_0_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_2_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o;
        end else begin
            l_TColl_0_2_1_constprop_o = l_TColl_0_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_2_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o;
        end else begin
            l_TColl_0_2_2_constprop_o = l_TColl_0_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_2_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o;
        end else begin
            l_TColl_0_2_3_constprop_o = l_TColl_0_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_3_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o;
        end else begin
            l_TColl_0_3_0_constprop_o = l_TColl_0_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_3_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o;
        end else begin
            l_TColl_0_3_1_constprop_o = l_TColl_0_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_3_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o;
        end else begin
            l_TColl_0_3_2_constprop_o = l_TColl_0_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_0_3_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o;
        end else begin
            l_TColl_0_3_3_constprop_o = l_TColl_0_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_0_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o;
        end else begin
            l_TColl_1_0_0_constprop_o = l_TColl_1_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_0_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o;
        end else begin
            l_TColl_1_0_1_constprop_o = l_TColl_1_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_0_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o;
        end else begin
            l_TColl_1_0_2_constprop_o = l_TColl_1_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_0_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o;
        end else begin
            l_TColl_1_0_3_constprop_o = l_TColl_1_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_1_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o;
        end else begin
            l_TColl_1_1_0_constprop_o = l_TColl_1_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_1_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o;
        end else begin
            l_TColl_1_1_1_constprop_o = l_TColl_1_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_1_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o;
        end else begin
            l_TColl_1_1_2_constprop_o = l_TColl_1_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_1_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o;
        end else begin
            l_TColl_1_1_3_constprop_o = l_TColl_1_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_2_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o;
        end else begin
            l_TColl_1_2_0_constprop_o = l_TColl_1_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_2_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o;
        end else begin
            l_TColl_1_2_1_constprop_o = l_TColl_1_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_2_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o;
        end else begin
            l_TColl_1_2_2_constprop_o = l_TColl_1_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_2_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o;
        end else begin
            l_TColl_1_2_3_constprop_o = l_TColl_1_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_3_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o;
        end else begin
            l_TColl_1_3_0_constprop_o = l_TColl_1_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_3_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o;
        end else begin
            l_TColl_1_3_1_constprop_o = l_TColl_1_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_3_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o;
        end else begin
            l_TColl_1_3_2_constprop_o = l_TColl_1_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_1_3_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o;
        end else begin
            l_TColl_1_3_3_constprop_o = l_TColl_1_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_0_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o;
        end else begin
            l_TColl_2_0_0_constprop_o = l_TColl_2_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_0_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o;
        end else begin
            l_TColl_2_0_1_constprop_o = l_TColl_2_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_0_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o;
        end else begin
            l_TColl_2_0_2_constprop_o = l_TColl_2_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_0_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o;
        end else begin
            l_TColl_2_0_3_constprop_o = l_TColl_2_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_1_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o;
        end else begin
            l_TColl_2_1_0_constprop_o = l_TColl_2_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_1_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o;
        end else begin
            l_TColl_2_1_1_constprop_o = l_TColl_2_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_1_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o;
        end else begin
            l_TColl_2_1_2_constprop_o = l_TColl_2_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_1_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o;
        end else begin
            l_TColl_2_1_3_constprop_o = l_TColl_2_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_2_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o;
        end else begin
            l_TColl_2_2_0_constprop_o = l_TColl_2_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_2_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o;
        end else begin
            l_TColl_2_2_1_constprop_o = l_TColl_2_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_2_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o;
        end else begin
            l_TColl_2_2_2_constprop_o = l_TColl_2_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_2_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o;
        end else begin
            l_TColl_2_2_3_constprop_o = l_TColl_2_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_3_0_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o;
        end else begin
            l_TColl_2_3_0_constprop_o = l_TColl_2_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_3_1_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o;
        end else begin
            l_TColl_2_3_1_constprop_o = l_TColl_2_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_3_2_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o;
        end else begin
            l_TColl_2_3_2_constprop_o = l_TColl_2_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o_ap_vld == 1'b1))) begin
            l_TColl_2_3_3_constprop_o = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o;
        end else begin
            l_TColl_2_3_3_constprop_o = l_TColl_2_3_3_constprop_i;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_0_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_0_address0 = grp_forwardKin_fu_863_this_TCurr_0_0_address0;
        end else begin
            this_TCurr_0_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_0_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_0_ce0 = grp_forwardKin_fu_863_this_TCurr_0_0_ce0;
        end else begin
            this_TCurr_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_0_we0 = grp_forwardKin_fu_863_this_TCurr_0_0_we0;
        end else begin
            this_TCurr_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_1_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_1_address0 = grp_forwardKin_fu_863_this_TCurr_0_1_address0;
        end else begin
            this_TCurr_0_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_1_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_1_ce0 = grp_forwardKin_fu_863_this_TCurr_0_1_ce0;
        end else begin
            this_TCurr_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_1_we0 = grp_forwardKin_fu_863_this_TCurr_0_1_we0;
        end else begin
            this_TCurr_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_2_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_2_address0 = grp_forwardKin_fu_863_this_TCurr_0_2_address0;
        end else begin
            this_TCurr_0_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_2_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_2_ce0 = grp_forwardKin_fu_863_this_TCurr_0_2_ce0;
        end else begin
            this_TCurr_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_2_we0 = grp_forwardKin_fu_863_this_TCurr_0_2_we0;
        end else begin
            this_TCurr_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_3_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_3_address0 = grp_forwardKin_fu_863_this_TCurr_0_3_address0;
        end else begin
            this_TCurr_0_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_0_3_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_0_3_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_3_ce0 = grp_forwardKin_fu_863_this_TCurr_0_3_ce0;
        end else begin
            this_TCurr_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_0_3_we0 = grp_forwardKin_fu_863_this_TCurr_0_3_we0;
        end else begin
            this_TCurr_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_0_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_0_address0 = grp_forwardKin_fu_863_this_TCurr_1_0_address0;
        end else begin
            this_TCurr_1_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_0_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_0_ce0 = grp_forwardKin_fu_863_this_TCurr_1_0_ce0;
        end else begin
            this_TCurr_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_0_we0 = grp_forwardKin_fu_863_this_TCurr_1_0_we0;
        end else begin
            this_TCurr_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_1_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_1_address0 = grp_forwardKin_fu_863_this_TCurr_1_1_address0;
        end else begin
            this_TCurr_1_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_1_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_1_ce0 = grp_forwardKin_fu_863_this_TCurr_1_1_ce0;
        end else begin
            this_TCurr_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_1_we0 = grp_forwardKin_fu_863_this_TCurr_1_1_we0;
        end else begin
            this_TCurr_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_2_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_2_address0 = grp_forwardKin_fu_863_this_TCurr_1_2_address0;
        end else begin
            this_TCurr_1_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_2_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_2_ce0 = grp_forwardKin_fu_863_this_TCurr_1_2_ce0;
        end else begin
            this_TCurr_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_2_we0 = grp_forwardKin_fu_863_this_TCurr_1_2_we0;
        end else begin
            this_TCurr_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_3_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_3_address0 = grp_forwardKin_fu_863_this_TCurr_1_3_address0;
        end else begin
            this_TCurr_1_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_1_3_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_1_3_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_3_ce0 = grp_forwardKin_fu_863_this_TCurr_1_3_ce0;
        end else begin
            this_TCurr_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_1_3_we0 = grp_forwardKin_fu_863_this_TCurr_1_3_we0;
        end else begin
            this_TCurr_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_0_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_0_address0 = grp_forwardKin_fu_863_this_TCurr_2_0_address0;
        end else begin
            this_TCurr_2_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_0_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_0_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_0_ce0 = grp_forwardKin_fu_863_this_TCurr_2_0_ce0;
        end else begin
            this_TCurr_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_0_we0 = grp_forwardKin_fu_863_this_TCurr_2_0_we0;
        end else begin
            this_TCurr_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_1_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_1_address0 = grp_forwardKin_fu_863_this_TCurr_2_1_address0;
        end else begin
            this_TCurr_2_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_1_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_1_ce0 = grp_forwardKin_fu_863_this_TCurr_2_1_ce0;
        end else begin
            this_TCurr_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_1_we0 = grp_forwardKin_fu_863_this_TCurr_2_1_we0;
        end else begin
            this_TCurr_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_2_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_2_address0 = grp_forwardKin_fu_863_this_TCurr_2_2_address0;
        end else begin
            this_TCurr_2_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_2_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_2_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_2_ce0 = grp_forwardKin_fu_863_this_TCurr_2_2_ce0;
        end else begin
            this_TCurr_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_2_we0 = grp_forwardKin_fu_863_this_TCurr_2_2_we0;
        end else begin
            this_TCurr_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_3_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_3_address0 = grp_forwardKin_fu_863_this_TCurr_2_3_address0;
        end else begin
            this_TCurr_2_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TCurr_2_3_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_TCurr_2_3_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_3_ce0 = grp_forwardKin_fu_863_this_TCurr_2_3_ce0;
        end else begin
            this_TCurr_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TCurr_2_3_we0 = grp_forwardKin_fu_863_this_TCurr_2_3_we0;
        end else begin
            this_TCurr_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cAxes_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cAxes_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_address0;
        end else begin
            this_cAxes_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cAxes_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cAxes_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_ce0;
        end else begin
            this_cAxes_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cAxes_ce1 = grp_cuboidCuboidCollision_double_s_fu_1252_axes1_ce1;
        end else begin
            this_cAxes_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cAxes_we0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_we0;
        end else begin
            this_cAxes_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cPoints_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p1_address0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_address0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address0;
        end else begin
            this_cPoints_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cPoints_address1 = grp_cuboidCuboidCollision_double_s_fu_1252_p1_address1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_address1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_address1;
        end else begin
            this_cPoints_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cPoints_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_ce0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce0;
        end else begin
            this_cPoints_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            this_cPoints_ce1 = grp_cuboidCuboidCollision_double_s_fu_1252_p1_ce1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_ce1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_ce1;
        end else begin
            this_cPoints_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_we0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we0;
        end else begin
            this_cPoints_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_cPoints_we1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_we1;
        end else begin
            this_cPoints_we1 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                if (((1'b1 == ap_CS_fsm_state2) & (1'b0 == ap_block_state2_on_subcall_done))) begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                if (((1'b1 == ap_CS_fsm_state4) & (grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            ap_ST_fsm_state5: begin
                if (((1'b1 == ap_CS_fsm_state5) & (icmp_ln168_fu_1327_p2 == 1'd0))) begin
                    ap_NS_fsm = ap_ST_fsm_state6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state8;
                end
            end
            ap_ST_fsm_state6: begin
                if (((1'b1 == ap_CS_fsm_state6) & (icmp_ln169_fu_1351_p2 == 1'd1))) begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state7;
                end
            end
            ap_ST_fsm_state7: begin
                if (((1'b1 == ap_CS_fsm_state7) & (grp_cuboidCuboidCollision_double_s_fu_1252_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state7;
                end
            end
            ap_ST_fsm_state8: begin
                if (((1'b1 == ap_CS_fsm_state8) & (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state8;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln168_fu_1333_p2 = (i_fu_448 + 3'd1);

    assign add_ln169_fu_1357_p2 = (j_reg_852 + 4'd1);

    assign add_ln170_fu_1372_p2 = (zext_ln169_fu_1363_p1 + tmp_48_reg_1731);

    assign ang_address0 = grp_forwardKin_fu_863_ang_address0;

    assign ang_ce0 = grp_forwardKin_fu_863_ang_ce0;

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    always @(*) begin
        ap_block_state2_on_subcall_done = ((grp_forwardKin_fu_863_ap_done == 1'b0) | (grp_detectCollNode_Pipeline_2_fu_985_ap_done == 1'b0));
    end

    assign grp_cuboidCuboidCollision_double_s_fu_1252_ap_start = grp_cuboidCuboidCollision_double_s_fu_1252_ap_start_reg;

    assign grp_detectCollNode_Pipeline_2_fu_985_ap_start = grp_detectCollNode_Pipeline_2_fu_985_ap_start_reg;

    assign grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start = grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_start_reg;

    assign grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_ap_start_reg;

    assign grp_forwardKin_fu_863_ap_start = grp_forwardKin_fu_863_ap_start_reg;

    assign grp_fu_1454_p_ce = grp_fu_1794_ce;

    assign grp_fu_1454_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din0;

    assign grp_fu_1454_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_din1;

    assign grp_fu_1454_p_opcode = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1794_p_opcode;

    assign grp_fu_1462_p_ce = grp_fu_1798_ce;

    assign grp_fu_1462_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din0;

    assign grp_fu_1462_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1798_p_din1;

    assign grp_fu_2529_p_ce = grp_fu_1754_ce;

    assign grp_fu_2529_p_din0 = grp_fu_1754_p0;

    assign grp_fu_2529_p_din1 = grp_fu_1754_p1;

    assign grp_fu_2529_p_opcode = grp_fu_1754_opcode;

    assign grp_fu_2533_p_ce = grp_fu_1758_ce;

    assign grp_fu_2533_p_din0 = grp_fu_1758_p0;

    assign grp_fu_2533_p_din1 = grp_fu_1758_p1;

    assign grp_fu_2537_p_ce = grp_fu_1762_ce;

    assign grp_fu_2537_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din0;

    assign grp_fu_2537_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_din1;

    assign grp_fu_2537_p_opcode = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1762_p_opcode;

    assign grp_fu_2541_p_ce = grp_fu_1766_ce;

    assign grp_fu_2541_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din0;

    assign grp_fu_2541_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_din1;

    assign grp_fu_2541_p_opcode = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1766_p_opcode;

    assign grp_fu_2545_p_ce = grp_fu_1770_ce;

    assign grp_fu_2545_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din0;

    assign grp_fu_2545_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1770_p_din1;

    assign grp_fu_2545_p_opcode = 2'd0;

    assign grp_fu_2549_p_ce = grp_fu_1774_ce;

    assign grp_fu_2549_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din0;

    assign grp_fu_2549_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1774_p_din1;

    assign grp_fu_2549_p_opcode = 2'd0;

    assign grp_fu_2553_p_ce = grp_fu_1778_ce;

    assign grp_fu_2553_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din0;

    assign grp_fu_2553_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1778_p_din1;

    assign grp_fu_2553_p_opcode = 2'd0;

    assign grp_fu_2557_p_ce = grp_fu_1782_ce;

    assign grp_fu_2557_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din0;

    assign grp_fu_2557_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1782_p_din1;

    assign grp_fu_2561_p_ce = grp_fu_1786_ce;

    assign grp_fu_2561_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din0;

    assign grp_fu_2561_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1786_p_din1;

    assign grp_fu_2565_p_ce = grp_fu_1790_ce;

    assign grp_fu_2565_p_din0 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din0;

    assign grp_fu_2565_p_din1 = grp_cuboidCuboidCollision_double_s_fu_1252_grp_fu_1790_p_din1;

    assign icmp_ln168_fu_1327_p2 = ((i_fu_448 == 3'd4) ? 1'b1 : 1'b0);

    assign icmp_ln169_fu_1351_p2 = ((j_reg_852 == 4'd8) ? 1'b1 : 1'b0);

    assign l_TColl_0_0_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_0_constprop_o_ap_vld;

    assign l_TColl_0_0_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_1_constprop_o_ap_vld;

    assign l_TColl_0_0_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_2_constprop_o_ap_vld;

    assign l_TColl_0_0_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_0_3_constprop_o_ap_vld;

    assign l_TColl_0_1_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_0_constprop_o_ap_vld;

    assign l_TColl_0_1_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_1_constprop_o_ap_vld;

    assign l_TColl_0_1_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_2_constprop_o_ap_vld;

    assign l_TColl_0_1_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_1_3_constprop_o_ap_vld;

    assign l_TColl_0_2_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_0_constprop_o_ap_vld;

    assign l_TColl_0_2_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_1_constprop_o_ap_vld;

    assign l_TColl_0_2_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_2_constprop_o_ap_vld;

    assign l_TColl_0_2_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_2_3_constprop_o_ap_vld;

    assign l_TColl_0_3_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_0_constprop_o_ap_vld;

    assign l_TColl_0_3_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_1_constprop_o_ap_vld;

    assign l_TColl_0_3_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_2_constprop_o_ap_vld;

    assign l_TColl_0_3_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_0_3_3_constprop_o_ap_vld;

    assign l_TColl_1_0_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_0_constprop_o_ap_vld;

    assign l_TColl_1_0_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_1_constprop_o_ap_vld;

    assign l_TColl_1_0_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_2_constprop_o_ap_vld;

    assign l_TColl_1_0_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_0_3_constprop_o_ap_vld;

    assign l_TColl_1_1_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_0_constprop_o_ap_vld;

    assign l_TColl_1_1_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_1_constprop_o_ap_vld;

    assign l_TColl_1_1_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_2_constprop_o_ap_vld;

    assign l_TColl_1_1_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_1_3_constprop_o_ap_vld;

    assign l_TColl_1_2_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_0_constprop_o_ap_vld;

    assign l_TColl_1_2_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_1_constprop_o_ap_vld;

    assign l_TColl_1_2_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_2_constprop_o_ap_vld;

    assign l_TColl_1_2_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_2_3_constprop_o_ap_vld;

    assign l_TColl_1_3_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_0_constprop_o_ap_vld;

    assign l_TColl_1_3_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_1_constprop_o_ap_vld;

    assign l_TColl_1_3_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_2_constprop_o_ap_vld;

    assign l_TColl_1_3_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_1_3_3_constprop_o_ap_vld;

    assign l_TColl_2_0_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_0_constprop_o_ap_vld;

    assign l_TColl_2_0_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_1_constprop_o_ap_vld;

    assign l_TColl_2_0_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_2_constprop_o_ap_vld;

    assign l_TColl_2_0_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_0_3_constprop_o_ap_vld;

    assign l_TColl_2_1_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_0_constprop_o_ap_vld;

    assign l_TColl_2_1_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_1_constprop_o_ap_vld;

    assign l_TColl_2_1_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_2_constprop_o_ap_vld;

    assign l_TColl_2_1_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_1_3_constprop_o_ap_vld;

    assign l_TColl_2_2_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_0_constprop_o_ap_vld;

    assign l_TColl_2_2_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_1_constprop_o_ap_vld;

    assign l_TColl_2_2_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_2_constprop_o_ap_vld;

    assign l_TColl_2_2_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_2_3_constprop_o_ap_vld;

    assign l_TColl_2_3_0_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_0_constprop_o_ap_vld;

    assign l_TColl_2_3_1_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_1_constprop_o_ap_vld;

    assign l_TColl_2_3_2_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_2_constprop_o_ap_vld;

    assign l_TColl_2_3_3_constprop_o_ap_vld = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_l_TColl_2_3_3_constprop_o_ap_vld;

    assign this_TCurr_0_0_d0 = grp_forwardKin_fu_863_this_TCurr_0_0_d0;

    assign this_TCurr_0_1_d0 = grp_forwardKin_fu_863_this_TCurr_0_1_d0;

    assign this_TCurr_0_2_d0 = grp_forwardKin_fu_863_this_TCurr_0_2_d0;

    assign this_TCurr_0_3_d0 = grp_forwardKin_fu_863_this_TCurr_0_3_d0;

    assign this_TCurr_1_0_d0 = grp_forwardKin_fu_863_this_TCurr_1_0_d0;

    assign this_TCurr_1_1_d0 = grp_forwardKin_fu_863_this_TCurr_1_1_d0;

    assign this_TCurr_1_2_d0 = grp_forwardKin_fu_863_this_TCurr_1_2_d0;

    assign this_TCurr_1_3_d0 = grp_forwardKin_fu_863_this_TCurr_1_3_d0;

    assign this_TCurr_2_0_d0 = grp_forwardKin_fu_863_this_TCurr_2_0_d0;

    assign this_TCurr_2_1_d0 = grp_forwardKin_fu_863_this_TCurr_2_1_d0;

    assign this_TCurr_2_2_d0 = grp_forwardKin_fu_863_this_TCurr_2_2_d0;

    assign this_TCurr_2_3_d0 = grp_forwardKin_fu_863_this_TCurr_2_3_d0;

    assign this_TCurr_3_0_address0 = grp_forwardKin_fu_863_this_TCurr_3_0_address0;

    assign this_TCurr_3_0_ce0 = grp_forwardKin_fu_863_this_TCurr_3_0_ce0;

    assign this_TCurr_3_0_d0 = grp_forwardKin_fu_863_this_TCurr_3_0_d0;

    assign this_TCurr_3_0_we0 = grp_forwardKin_fu_863_this_TCurr_3_0_we0;

    assign this_TCurr_3_1_address0 = grp_forwardKin_fu_863_this_TCurr_3_1_address0;

    assign this_TCurr_3_1_ce0 = grp_forwardKin_fu_863_this_TCurr_3_1_ce0;

    assign this_TCurr_3_1_d0 = grp_forwardKin_fu_863_this_TCurr_3_1_d0;

    assign this_TCurr_3_1_we0 = grp_forwardKin_fu_863_this_TCurr_3_1_we0;

    assign this_TCurr_3_2_address0 = grp_forwardKin_fu_863_this_TCurr_3_2_address0;

    assign this_TCurr_3_2_ce0 = grp_forwardKin_fu_863_this_TCurr_3_2_ce0;

    assign this_TCurr_3_2_d0 = grp_forwardKin_fu_863_this_TCurr_3_2_d0;

    assign this_TCurr_3_2_we0 = grp_forwardKin_fu_863_this_TCurr_3_2_we0;

    assign this_TCurr_3_3_address0 = grp_forwardKin_fu_863_this_TCurr_3_3_address0;

    assign this_TCurr_3_3_ce0 = grp_forwardKin_fu_863_this_TCurr_3_3_ce0;

    assign this_TCurr_3_3_d0 = grp_forwardKin_fu_863_this_TCurr_3_3_d0;

    assign this_TCurr_3_3_we0 = grp_forwardKin_fu_863_this_TCurr_3_3_we0;

    assign this_TJoint_0_0_address0 = grp_forwardKin_fu_863_this_TJoint_0_0_address0;

    assign this_TJoint_0_0_ce0 = grp_forwardKin_fu_863_this_TJoint_0_0_ce0;

    assign this_TJoint_0_0_d0 = grp_forwardKin_fu_863_this_TJoint_0_0_d0;

    assign this_TJoint_0_0_we0 = grp_forwardKin_fu_863_this_TJoint_0_0_we0;

    assign this_TJoint_0_1_address0 = grp_forwardKin_fu_863_this_TJoint_0_1_address0;

    assign this_TJoint_0_1_ce0 = grp_forwardKin_fu_863_this_TJoint_0_1_ce0;

    assign this_TJoint_0_1_d0 = grp_forwardKin_fu_863_this_TJoint_0_1_d0;

    assign this_TJoint_0_1_we0 = grp_forwardKin_fu_863_this_TJoint_0_1_we0;

    assign this_TJoint_0_2_address0 = grp_forwardKin_fu_863_this_TJoint_0_2_address0;

    assign this_TJoint_0_2_ce0 = grp_forwardKin_fu_863_this_TJoint_0_2_ce0;

    assign this_TJoint_0_2_d0 = grp_forwardKin_fu_863_this_TJoint_0_2_d0;

    assign this_TJoint_0_2_we0 = grp_forwardKin_fu_863_this_TJoint_0_2_we0;

    assign this_TJoint_0_3_address0 = grp_forwardKin_fu_863_this_TJoint_0_3_address0;

    assign this_TJoint_0_3_ce0 = grp_forwardKin_fu_863_this_TJoint_0_3_ce0;

    assign this_TJoint_0_3_d0 = grp_forwardKin_fu_863_this_TJoint_0_3_d0;

    assign this_TJoint_0_3_we0 = grp_forwardKin_fu_863_this_TJoint_0_3_we0;

    assign this_TJoint_1_0_address0 = grp_forwardKin_fu_863_this_TJoint_1_0_address0;

    assign this_TJoint_1_0_ce0 = grp_forwardKin_fu_863_this_TJoint_1_0_ce0;

    assign this_TJoint_1_0_d0 = grp_forwardKin_fu_863_this_TJoint_1_0_d0;

    assign this_TJoint_1_0_we0 = grp_forwardKin_fu_863_this_TJoint_1_0_we0;

    assign this_TJoint_1_1_address0 = grp_forwardKin_fu_863_this_TJoint_1_1_address0;

    assign this_TJoint_1_1_ce0 = grp_forwardKin_fu_863_this_TJoint_1_1_ce0;

    assign this_TJoint_1_1_d0 = grp_forwardKin_fu_863_this_TJoint_1_1_d0;

    assign this_TJoint_1_1_we0 = grp_forwardKin_fu_863_this_TJoint_1_1_we0;

    assign this_TJoint_1_2_address0 = grp_forwardKin_fu_863_this_TJoint_1_2_address0;

    assign this_TJoint_1_2_ce0 = grp_forwardKin_fu_863_this_TJoint_1_2_ce0;

    assign this_TJoint_1_2_d0 = grp_forwardKin_fu_863_this_TJoint_1_2_d0;

    assign this_TJoint_1_2_we0 = grp_forwardKin_fu_863_this_TJoint_1_2_we0;

    assign this_TJoint_1_3_address0 = grp_forwardKin_fu_863_this_TJoint_1_3_address0;

    assign this_TJoint_1_3_ce0 = grp_forwardKin_fu_863_this_TJoint_1_3_ce0;

    assign this_TJoint_1_3_d0 = grp_forwardKin_fu_863_this_TJoint_1_3_d0;

    assign this_TJoint_1_3_we0 = grp_forwardKin_fu_863_this_TJoint_1_3_we0;

    assign this_TJoint_2_0_address0 = grp_forwardKin_fu_863_this_TJoint_2_0_address0;

    assign this_TJoint_2_0_ce0 = grp_forwardKin_fu_863_this_TJoint_2_0_ce0;

    assign this_TJoint_2_0_d0 = grp_forwardKin_fu_863_this_TJoint_2_0_d0;

    assign this_TJoint_2_0_we0 = grp_forwardKin_fu_863_this_TJoint_2_0_we0;

    assign this_TJoint_2_1_address0 = grp_forwardKin_fu_863_this_TJoint_2_1_address0;

    assign this_TJoint_2_1_ce0 = grp_forwardKin_fu_863_this_TJoint_2_1_ce0;

    assign this_TJoint_2_1_d0 = grp_forwardKin_fu_863_this_TJoint_2_1_d0;

    assign this_TJoint_2_1_we0 = grp_forwardKin_fu_863_this_TJoint_2_1_we0;

    assign this_TJoint_2_2_address0 = grp_forwardKin_fu_863_this_TJoint_2_2_address0;

    assign this_TJoint_2_2_ce0 = grp_forwardKin_fu_863_this_TJoint_2_2_ce0;

    assign this_TJoint_2_2_d0 = grp_forwardKin_fu_863_this_TJoint_2_2_d0;

    assign this_TJoint_2_2_we0 = grp_forwardKin_fu_863_this_TJoint_2_2_we0;

    assign this_TJoint_2_3_address0 = grp_forwardKin_fu_863_this_TJoint_2_3_address0;

    assign this_TJoint_2_3_ce0 = grp_forwardKin_fu_863_this_TJoint_2_3_ce0;

    assign this_TJoint_2_3_d0 = grp_forwardKin_fu_863_this_TJoint_2_3_d0;

    assign this_TJoint_2_3_we0 = grp_forwardKin_fu_863_this_TJoint_2_3_we0;

    assign this_TJoint_3_0_address0 = grp_forwardKin_fu_863_this_TJoint_3_0_address0;

    assign this_TJoint_3_0_ce0 = grp_forwardKin_fu_863_this_TJoint_3_0_ce0;

    assign this_TJoint_3_0_d0 = grp_forwardKin_fu_863_this_TJoint_3_0_d0;

    assign this_TJoint_3_0_we0 = grp_forwardKin_fu_863_this_TJoint_3_0_we0;

    assign this_TJoint_3_1_address0 = grp_forwardKin_fu_863_this_TJoint_3_1_address0;

    assign this_TJoint_3_1_ce0 = grp_forwardKin_fu_863_this_TJoint_3_1_ce0;

    assign this_TJoint_3_1_d0 = grp_forwardKin_fu_863_this_TJoint_3_1_d0;

    assign this_TJoint_3_1_we0 = grp_forwardKin_fu_863_this_TJoint_3_1_we0;

    assign this_TJoint_3_2_address0 = grp_forwardKin_fu_863_this_TJoint_3_2_address0;

    assign this_TJoint_3_2_ce0 = grp_forwardKin_fu_863_this_TJoint_3_2_ce0;

    assign this_TJoint_3_2_d0 = grp_forwardKin_fu_863_this_TJoint_3_2_d0;

    assign this_TJoint_3_2_we0 = grp_forwardKin_fu_863_this_TJoint_3_2_we0;

    assign this_TJoint_3_3_address0 = grp_forwardKin_fu_863_this_TJoint_3_3_address0;

    assign this_TJoint_3_3_ce0 = grp_forwardKin_fu_863_this_TJoint_3_3_ce0;

    assign this_TJoint_3_3_d0 = grp_forwardKin_fu_863_this_TJoint_3_3_d0;

    assign this_TJoint_3_3_we0 = grp_forwardKin_fu_863_this_TJoint_3_3_we0;

    assign this_TLink_0_0_address0 = grp_forwardKin_fu_863_this_TLink_0_0_address0;

    assign this_TLink_0_0_ce0 = grp_forwardKin_fu_863_this_TLink_0_0_ce0;

    assign this_TLink_0_1_address0 = grp_forwardKin_fu_863_this_TLink_0_1_address0;

    assign this_TLink_0_1_ce0 = grp_forwardKin_fu_863_this_TLink_0_1_ce0;

    assign this_TLink_0_2_address0 = grp_forwardKin_fu_863_this_TLink_0_2_address0;

    assign this_TLink_0_2_ce0 = grp_forwardKin_fu_863_this_TLink_0_2_ce0;

    assign this_TLink_0_3_address0 = grp_forwardKin_fu_863_this_TLink_0_3_address0;

    assign this_TLink_0_3_ce0 = grp_forwardKin_fu_863_this_TLink_0_3_ce0;

    assign this_TLink_1_0_address0 = grp_forwardKin_fu_863_this_TLink_1_0_address0;

    assign this_TLink_1_0_ce0 = grp_forwardKin_fu_863_this_TLink_1_0_ce0;

    assign this_TLink_1_1_address0 = grp_forwardKin_fu_863_this_TLink_1_1_address0;

    assign this_TLink_1_1_ce0 = grp_forwardKin_fu_863_this_TLink_1_1_ce0;

    assign this_TLink_1_2_address0 = grp_forwardKin_fu_863_this_TLink_1_2_address0;

    assign this_TLink_1_2_ce0 = grp_forwardKin_fu_863_this_TLink_1_2_ce0;

    assign this_TLink_1_3_address0 = grp_forwardKin_fu_863_this_TLink_1_3_address0;

    assign this_TLink_1_3_ce0 = grp_forwardKin_fu_863_this_TLink_1_3_ce0;

    assign this_TLink_2_0_address0 = grp_forwardKin_fu_863_this_TLink_2_0_address0;

    assign this_TLink_2_0_ce0 = grp_forwardKin_fu_863_this_TLink_2_0_ce0;

    assign this_TLink_2_1_address0 = grp_forwardKin_fu_863_this_TLink_2_1_address0;

    assign this_TLink_2_1_ce0 = grp_forwardKin_fu_863_this_TLink_2_1_ce0;

    assign this_TLink_2_2_address0 = grp_forwardKin_fu_863_this_TLink_2_2_address0;

    assign this_TLink_2_2_ce0 = grp_forwardKin_fu_863_this_TLink_2_2_ce0;

    assign this_TLink_2_3_address0 = grp_forwardKin_fu_863_this_TLink_2_3_address0;

    assign this_TLink_2_3_ce0 = grp_forwardKin_fu_863_this_TLink_2_3_ce0;

    assign this_TLink_3_0_address0 = grp_forwardKin_fu_863_this_TLink_3_0_address0;

    assign this_TLink_3_0_ce0 = grp_forwardKin_fu_863_this_TLink_3_0_ce0;

    assign this_TLink_3_1_address0 = grp_forwardKin_fu_863_this_TLink_3_1_address0;

    assign this_TLink_3_1_ce0 = grp_forwardKin_fu_863_this_TLink_3_1_ce0;

    assign this_TLink_3_2_address0 = grp_forwardKin_fu_863_this_TLink_3_2_address0;

    assign this_TLink_3_2_ce0 = grp_forwardKin_fu_863_this_TLink_3_2_ce0;

    assign this_TLink_3_3_address0 = grp_forwardKin_fu_863_this_TLink_3_3_address0;

    assign this_TLink_3_3_ce0 = grp_forwardKin_fu_863_this_TLink_3_3_ce0;

    assign this_cAxes_address1 = grp_cuboidCuboidCollision_double_s_fu_1252_axes1_address1;

    assign this_cAxes_d0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cAxes_d0;

    assign this_cPoints_d0 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d0;

    assign this_cPoints_d1 = grp_detectCollNode_Pipeline_VITIS_LOOP_276_1_fu_991_this_cPoints_d1;

    assign this_env_0_0_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_address0;

    assign this_env_0_0_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_0_ce0;

    assign this_env_0_0_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_address0;

    assign this_env_0_0_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_1_ce0;

    assign this_env_0_0_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_address0;

    assign this_env_0_0_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_0_2_ce0;

    assign this_env_0_1_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_address0;

    assign this_env_0_1_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_0_ce0;

    assign this_env_0_1_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_address0;

    assign this_env_0_1_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_1_ce0;

    assign this_env_0_1_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_address0;

    assign this_env_0_1_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_1_2_ce0;

    assign this_env_0_2_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_address0;

    assign this_env_0_2_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_0_ce0;

    assign this_env_0_2_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_address0;

    assign this_env_0_2_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_1_ce0;

    assign this_env_0_2_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_address0;

    assign this_env_0_2_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_2_2_ce0;

    assign this_env_0_3_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_address0;

    assign this_env_0_3_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_0_ce0;

    assign this_env_0_3_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_address0;

    assign this_env_0_3_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_1_ce0;

    assign this_env_0_3_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_address0;

    assign this_env_0_3_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_3_2_ce0;

    assign this_env_0_4_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_address0;

    assign this_env_0_4_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_0_ce0;

    assign this_env_0_4_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_address0;

    assign this_env_0_4_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_1_ce0;

    assign this_env_0_4_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_address0;

    assign this_env_0_4_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_4_2_ce0;

    assign this_env_0_5_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_address0;

    assign this_env_0_5_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_0_ce0;

    assign this_env_0_5_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_address0;

    assign this_env_0_5_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_1_ce0;

    assign this_env_0_5_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_address0;

    assign this_env_0_5_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_5_2_ce0;

    assign this_env_0_6_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_address0;

    assign this_env_0_6_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_0_ce0;

    assign this_env_0_6_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_address0;

    assign this_env_0_6_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_1_ce0;

    assign this_env_0_6_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_address0;

    assign this_env_0_6_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_6_2_ce0;

    assign this_env_0_7_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_address0;

    assign this_env_0_7_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_0_ce0;

    assign this_env_0_7_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_address0;

    assign this_env_0_7_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_1_ce0;

    assign this_env_0_7_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_address0;

    assign this_env_0_7_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_7_2_ce0;

    assign this_env_0_8_0_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_address0;

    assign this_env_0_8_0_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_0_ce0;

    assign this_env_0_8_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_address0;

    assign this_env_0_8_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_1_ce0;

    assign this_env_0_8_2_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_address0;

    assign this_env_0_8_2_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_p2_8_2_ce0;

    assign this_env_1_address0 = grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address0;

    assign this_env_1_address1 = grp_cuboidCuboidCollision_double_s_fu_1252_axes2_address1;

    assign this_env_1_ce0 = grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce0;

    assign this_env_1_ce1 = grp_cuboidCuboidCollision_double_s_fu_1252_axes2_ce1;

    assign this_q_address0 = grp_forwardKin_fu_863_this_q_address0;

    assign this_q_ce0 = grp_forwardKin_fu_863_this_q_ce0;

    assign this_q_d0 = grp_forwardKin_fu_863_this_q_d0;

    assign this_q_we0 = grp_forwardKin_fu_863_this_q_we0;

    assign tmp_48_fu_1343_p3 = {{trunc_ln168_fu_1339_p1}, {3'd0}};

    assign trunc_ln168_fu_1339_p1 = i_fu_448[1:0];

    assign trunc_ln169_fu_1367_p1 = j_reg_852[2:0];

    assign xor_ln176_fu_1385_p2 = (grp_detectCollNode_Pipeline_VITIS_LOOP_176_3_fu_1247_ap_return ^ 1'd1);

    assign zext_ln169_fu_1363_p1 = j_reg_852;

    assign zext_ln170_fu_1381_p1 = add_ln170_reg_1749;

    always @(posedge ap_clk) begin
        tmp_48_reg_1731[2:0] <= 3'b000;
    end

endmodule  //main_detectCollNode
