/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    empty,
    axes1_address0,
    axes1_ce0,
    axes1_q0,
    axes1_address1,
    axes1_ce1,
    axes1_q1,
    sub_ln179,
    axes2_address0,
    axes2_ce0,
    axes2_q0,
    axes2_address1,
    axes2_ce1,
    axes2_q1,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    ap_return,
    grp_fu_469_p_din0,
    grp_fu_469_p_din1,
    grp_fu_469_p_opcode,
    grp_fu_469_p_dout0,
    grp_fu_469_p_ce,
    grp_fu_473_p_din0,
    grp_fu_473_p_din1,
    grp_fu_473_p_opcode,
    grp_fu_473_p_dout0,
    grp_fu_473_p_ce,
    grp_fu_493_p_din0,
    grp_fu_493_p_din1,
    grp_fu_493_p_dout0,
    grp_fu_493_p_ce,
    grp_fu_497_p_din0,
    grp_fu_497_p_din1,
    grp_fu_497_p_dout0,
    grp_fu_497_p_ce,
    grp_fu_501_p_din0,
    grp_fu_501_p_din1,
    grp_fu_501_p_dout0,
    grp_fu_501_p_ce,
    grp_fu_505_p_din0,
    grp_fu_505_p_din1,
    grp_fu_505_p_dout0,
    grp_fu_505_p_ce
);

    parameter ap_ST_fsm_state1 = 77'd1;
    parameter ap_ST_fsm_state2 = 77'd2;
    parameter ap_ST_fsm_state3 = 77'd4;
    parameter ap_ST_fsm_state4 = 77'd8;
    parameter ap_ST_fsm_state5 = 77'd16;
    parameter ap_ST_fsm_state6 = 77'd32;
    parameter ap_ST_fsm_state7 = 77'd64;
    parameter ap_ST_fsm_state8 = 77'd128;
    parameter ap_ST_fsm_state9 = 77'd256;
    parameter ap_ST_fsm_state10 = 77'd512;
    parameter ap_ST_fsm_state11 = 77'd1024;
    parameter ap_ST_fsm_state12 = 77'd2048;
    parameter ap_ST_fsm_state13 = 77'd4096;
    parameter ap_ST_fsm_state14 = 77'd8192;
    parameter ap_ST_fsm_state15 = 77'd16384;
    parameter ap_ST_fsm_state16 = 77'd32768;
    parameter ap_ST_fsm_state17 = 77'd65536;
    parameter ap_ST_fsm_state18 = 77'd131072;
    parameter ap_ST_fsm_state19 = 77'd262144;
    parameter ap_ST_fsm_state20 = 77'd524288;
    parameter ap_ST_fsm_state21 = 77'd1048576;
    parameter ap_ST_fsm_state22 = 77'd2097152;
    parameter ap_ST_fsm_state23 = 77'd4194304;
    parameter ap_ST_fsm_state24 = 77'd8388608;
    parameter ap_ST_fsm_state25 = 77'd16777216;
    parameter ap_ST_fsm_state26 = 77'd33554432;
    parameter ap_ST_fsm_state27 = 77'd67108864;
    parameter ap_ST_fsm_state28 = 77'd134217728;
    parameter ap_ST_fsm_state29 = 77'd268435456;
    parameter ap_ST_fsm_state30 = 77'd536870912;
    parameter ap_ST_fsm_state31 = 77'd1073741824;
    parameter ap_ST_fsm_state32 = 77'd2147483648;
    parameter ap_ST_fsm_state33 = 77'd4294967296;
    parameter ap_ST_fsm_state34 = 77'd8589934592;
    parameter ap_ST_fsm_state35 = 77'd17179869184;
    parameter ap_ST_fsm_state36 = 77'd34359738368;
    parameter ap_ST_fsm_state37 = 77'd68719476736;
    parameter ap_ST_fsm_state38 = 77'd137438953472;
    parameter ap_ST_fsm_state39 = 77'd274877906944;
    parameter ap_ST_fsm_state40 = 77'd549755813888;
    parameter ap_ST_fsm_state41 = 77'd1099511627776;
    parameter ap_ST_fsm_state42 = 77'd2199023255552;
    parameter ap_ST_fsm_state43 = 77'd4398046511104;
    parameter ap_ST_fsm_state44 = 77'd8796093022208;
    parameter ap_ST_fsm_state45 = 77'd17592186044416;
    parameter ap_ST_fsm_state46 = 77'd35184372088832;
    parameter ap_ST_fsm_state47 = 77'd70368744177664;
    parameter ap_ST_fsm_state48 = 77'd140737488355328;
    parameter ap_ST_fsm_state49 = 77'd281474976710656;
    parameter ap_ST_fsm_state50 = 77'd562949953421312;
    parameter ap_ST_fsm_state51 = 77'd1125899906842624;
    parameter ap_ST_fsm_state52 = 77'd2251799813685248;
    parameter ap_ST_fsm_state53 = 77'd4503599627370496;
    parameter ap_ST_fsm_state54 = 77'd9007199254740992;
    parameter ap_ST_fsm_state55 = 77'd18014398509481984;
    parameter ap_ST_fsm_state56 = 77'd36028797018963968;
    parameter ap_ST_fsm_state57 = 77'd72057594037927936;
    parameter ap_ST_fsm_state58 = 77'd144115188075855872;
    parameter ap_ST_fsm_state59 = 77'd288230376151711744;
    parameter ap_ST_fsm_state60 = 77'd576460752303423488;
    parameter ap_ST_fsm_state61 = 77'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 77'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 77'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 77'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 77'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 77'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 77'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 77'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 77'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 77'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 77'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 77'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 77'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 77'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 77'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 77'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 77'd75557863725914323419136;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [4:0] empty;
    output [5:0] axes1_address0;
    output axes1_ce0;
    input [63:0] axes1_q0;
    output [5:0] axes1_address1;
    output axes1_ce1;
    input [63:0] axes1_q1;
    input [5:0] sub_ln179;
    output [6:0] axes2_address0;
    output axes2_ce0;
    input [63:0] axes2_q0;
    output [6:0] axes2_address1;
    output axes2_ce1;
    input [63:0] axes2_q1;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    output [0:0] ap_return;
    output [63:0] grp_fu_469_p_din0;
    output [63:0] grp_fu_469_p_din1;
    output [0:0] grp_fu_469_p_opcode;
    input [63:0] grp_fu_469_p_dout0;
    output grp_fu_469_p_ce;
    output [63:0] grp_fu_473_p_din0;
    output [63:0] grp_fu_473_p_din1;
    output [0:0] grp_fu_473_p_opcode;
    input [63:0] grp_fu_473_p_dout0;
    output grp_fu_473_p_ce;
    output [63:0] grp_fu_493_p_din0;
    output [63:0] grp_fu_493_p_din1;
    input [63:0] grp_fu_493_p_dout0;
    output grp_fu_493_p_ce;
    output [63:0] grp_fu_497_p_din0;
    output [63:0] grp_fu_497_p_din1;
    input [63:0] grp_fu_497_p_dout0;
    output grp_fu_497_p_ce;
    output [63:0] grp_fu_501_p_din0;
    output [63:0] grp_fu_501_p_din1;
    input [63:0] grp_fu_501_p_dout0;
    output grp_fu_501_p_ce;
    output [63:0] grp_fu_505_p_din0;
    output [63:0] grp_fu_505_p_din1;
    input [63:0] grp_fu_505_p_dout0;
    output grp_fu_505_p_ce;

    reg ap_idle;
    reg[5:0] axes1_address0;
    reg axes1_ce0;
    reg axes1_ce1;
    reg[6:0] axes2_address0;
    reg axes2_ce0;
    reg axes2_ce1;
    reg[0:0] ap_return;

    (* fsm_encoding = "none" *) reg   [76:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire    ap_CS_fsm_state77;
    wire   [0:0] grp_pointsOverlap_double_s_fu_238_ap_return;
    reg   [0:0] icmp_ln184_reg_573;
    reg    ap_condition_exit_pp0_iter0_stage76;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    reg   [0:0] merge_reg_226;
    reg    ap_block_state1_pp0_stage0_iter0;
    reg   [1:0] i_reg_568;
    wire   [0:0] icmp_ln184_fu_378_p2;
    wire   [3:0] add_ln184_3_fu_384_p2;
    reg   [3:0] add_ln184_3_reg_577;
    wire   [1:0] add_ln184_fu_393_p2;
    reg   [1:0] add_ln184_reg_582;
    wire   [0:0] icmp_ln185_fu_399_p2;
    reg   [0:0] icmp_ln185_reg_587;
    wire   [1:0] select_ln184_fu_405_p3;
    reg   [1:0] select_ln184_reg_592;
    wire   [5:0] select_ln184_1_fu_435_p3;
    reg   [5:0] select_ln184_1_reg_597;
    wire   [6:0] add_ln179_fu_447_p2;
    reg   [6:0] add_ln179_reg_604;
    wire    ap_CS_fsm_state2;
    wire   [6:0] sub_ln179_1_fu_478_p2;
    reg   [6:0] sub_ln179_1_reg_620;
    reg   [63:0] axes1_load_reg_635;
    wire    ap_CS_fsm_state3;
    reg   [63:0] axes1_load_1_reg_641;
    reg   [63:0] axes2_load_reg_657;
    reg   [63:0] axes2_load_1_reg_663;
    reg   [63:0] axes1_load_2_reg_669;
    wire    ap_CS_fsm_state4;
    reg   [63:0] axes2_load_2_reg_675;
    reg   [63:0] mul_i_reg_681;
    wire    ap_CS_fsm_state10;
    reg   [63:0] mul5_i_reg_686;
    reg   [63:0] mul9_i_reg_691;
    wire    ap_CS_fsm_state11;
    reg   [63:0] mul12_i_reg_696;
    reg   [63:0] mul17_i_reg_701;
    reg   [63:0] mul20_i_reg_706;
    reg   [63:0] cm_0_reg_711;
    wire    ap_CS_fsm_state17;
    reg   [63:0] cm_1_reg_716;
    wire    ap_CS_fsm_state18;
    reg   [63:0] cm_2_reg_721;
    wire    grp_pointsOverlap_double_s_fu_238_ap_start;
    wire    grp_pointsOverlap_double_s_fu_238_ap_done;
    wire    grp_pointsOverlap_double_s_fu_238_ap_idle;
    wire    grp_pointsOverlap_double_s_fu_238_ap_ready;
    wire   [6:0] grp_pointsOverlap_double_s_fu_238_p1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p1_ce0;
    wire   [6:0] grp_pointsOverlap_double_s_fu_238_p1_address1;
    wire    grp_pointsOverlap_double_s_fu_238_p1_ce1;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_0_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_0_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_0_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_0_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_0_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_0_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_1_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_1_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_1_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_1_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_1_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_1_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_2_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_2_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_2_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_2_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_2_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_2_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_3_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_3_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_3_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_3_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_3_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_3_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_4_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_4_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_4_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_4_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_4_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_4_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_5_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_5_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_5_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_5_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_5_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_5_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_6_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_6_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_6_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_6_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_6_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_6_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_7_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_7_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_7_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_7_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_7_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_7_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_8_0_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_8_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_8_1_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_8_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_s_fu_238_p2_8_2_address0;
    wire    grp_pointsOverlap_double_s_fu_238_p2_8_2_ce0;
    reg   [0:0] ap_phi_mux_merge_phi_fu_230_p4;
    reg    grp_pointsOverlap_double_s_fu_238_ap_start_reg;
    reg   [76:0] ap_NS_fsm;
    wire    ap_NS_fsm_state19;
    wire    ap_CS_fsm_state19;
    wire    ap_CS_fsm_state20;
    wire    ap_CS_fsm_state21;
    wire    ap_CS_fsm_state22;
    wire    ap_CS_fsm_state23;
    wire    ap_CS_fsm_state24;
    wire    ap_CS_fsm_state25;
    wire    ap_CS_fsm_state26;
    wire    ap_CS_fsm_state27;
    wire    ap_CS_fsm_state28;
    wire    ap_CS_fsm_state29;
    wire    ap_CS_fsm_state30;
    wire    ap_CS_fsm_state31;
    wire    ap_CS_fsm_state32;
    wire    ap_CS_fsm_state33;
    wire   [63:0] add_ln184_1_cast_fu_458_p1;
    wire   [63:0] add_ln184_2_cast_fu_468_p1;
    wire   [63:0] zext_ln179_2_fu_489_p1;
    wire   [63:0] zext_ln179_3_fu_500_p1;
    wire   [63:0] zext_ln184_fu_505_p1;
    wire   [63:0] zext_ln179_1_fu_509_p1;
    reg   [1:0] j_fu_124;
    wire   [1:0] add_ln185_fu_518_p2;
    wire    ap_loop_init;
    reg   [1:0] ap_sig_allocacmp_j_load;
    reg   [1:0] i_3_fu_128;
    wire   [1:0] select_ln184_2_fu_513_p3;
    reg   [1:0] ap_sig_allocacmp_i;
    reg   [3:0] indvar_flatten_fu_132;
    reg   [3:0] ap_sig_allocacmp_indvar_flatten_load;
    reg   [63:0] grp_fu_303_p0;
    reg   [63:0] grp_fu_303_p1;
    wire    ap_CS_fsm_state12;
    reg   [63:0] grp_fu_311_p0;
    reg   [63:0] grp_fu_311_p1;
    wire    ap_CS_fsm_state5;
    reg   [63:0] grp_fu_315_p0;
    reg   [63:0] grp_fu_315_p1;
    wire  signed [5:0] p_cast_fu_331_p1;
    wire   [5:0] i_3_cast_fu_356_p1;
    wire   [5:0] empty_80_fu_360_p2;
    wire   [5:0] empty_81_fu_366_p2;
    wire   [5:0] add_ln184_cast_fu_413_p1;
    wire   [5:0] empty_83_fu_417_p2;
    wire   [5:0] empty_84_fu_423_p2;
    wire   [5:0] empty_85_fu_429_p2;
    wire   [5:0] empty_82_fu_372_p2;
    wire  signed [6:0] sub_ln179_cast_fu_327_p1;
    wire   [6:0] zext_ln179_fu_443_p1;
    wire   [5:0] add_ln184_1_fu_453_p2;
    wire   [5:0] add_ln184_2_fu_463_p2;
    wire   [6:0] shl_ln179_fu_473_p2;
    wire   [6:0] add_ln179_1_fu_483_p2;
    wire   [6:0] add_ln179_2_fu_494_p2;
    reg   [0:0] ap_return_preg;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_ST_fsm_state62_blk;
    wire    ap_ST_fsm_state63_blk;
    wire    ap_ST_fsm_state64_blk;
    wire    ap_ST_fsm_state65_blk;
    wire    ap_ST_fsm_state66_blk;
    wire    ap_ST_fsm_state67_blk;
    wire    ap_ST_fsm_state68_blk;
    wire    ap_ST_fsm_state69_blk;
    wire    ap_ST_fsm_state70_blk;
    wire    ap_ST_fsm_state71_blk;
    wire    ap_ST_fsm_state72_blk;
    wire    ap_ST_fsm_state73_blk;
    wire    ap_ST_fsm_state74_blk;
    wire    ap_ST_fsm_state75_blk;
    wire    ap_ST_fsm_state76_blk;
    wire    ap_ST_fsm_state77_blk;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 77'd1;
        #0 grp_pointsOverlap_double_s_fu_238_ap_start_reg = 1'b0;
        #0 j_fu_124 = 2'd0;
        #0 i_3_fu_128 = 2'd0;
        #0 indvar_flatten_fu_132 = 4'd0;
        #0 ap_return_preg = 1'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_pointsOverlap_double_s grp_pointsOverlap_double_s_fu_238 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_pointsOverlap_double_s_fu_238_ap_start),
        .ap_done(grp_pointsOverlap_double_s_fu_238_ap_done),
        .ap_idle(grp_pointsOverlap_double_s_fu_238_ap_idle),
        .ap_ready(grp_pointsOverlap_double_s_fu_238_ap_ready),
        .p1_address0(grp_pointsOverlap_double_s_fu_238_p1_address0),
        .p1_ce0(grp_pointsOverlap_double_s_fu_238_p1_ce0),
        .p1_q0(p1_q0),
        .p1_address1(grp_pointsOverlap_double_s_fu_238_p1_address1),
        .p1_ce1(grp_pointsOverlap_double_s_fu_238_p1_ce1),
        .p1_q1(p1_q1),
        .p1_offset(p1_offset),
        .p2_0_0_address0(grp_pointsOverlap_double_s_fu_238_p2_0_0_address0),
        .p2_0_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_0_0_ce0),
        .p2_0_0_q0(p2_0_0_q0),
        .p2_0_1_address0(grp_pointsOverlap_double_s_fu_238_p2_0_1_address0),
        .p2_0_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_0_1_ce0),
        .p2_0_1_q0(p2_0_1_q0),
        .p2_0_2_address0(grp_pointsOverlap_double_s_fu_238_p2_0_2_address0),
        .p2_0_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_0_2_ce0),
        .p2_0_2_q0(p2_0_2_q0),
        .p2_1_0_address0(grp_pointsOverlap_double_s_fu_238_p2_1_0_address0),
        .p2_1_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_1_0_ce0),
        .p2_1_0_q0(p2_1_0_q0),
        .p2_1_1_address0(grp_pointsOverlap_double_s_fu_238_p2_1_1_address0),
        .p2_1_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_1_1_ce0),
        .p2_1_1_q0(p2_1_1_q0),
        .p2_1_2_address0(grp_pointsOverlap_double_s_fu_238_p2_1_2_address0),
        .p2_1_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_1_2_ce0),
        .p2_1_2_q0(p2_1_2_q0),
        .p2_2_0_address0(grp_pointsOverlap_double_s_fu_238_p2_2_0_address0),
        .p2_2_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_2_0_ce0),
        .p2_2_0_q0(p2_2_0_q0),
        .p2_2_1_address0(grp_pointsOverlap_double_s_fu_238_p2_2_1_address0),
        .p2_2_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_2_1_ce0),
        .p2_2_1_q0(p2_2_1_q0),
        .p2_2_2_address0(grp_pointsOverlap_double_s_fu_238_p2_2_2_address0),
        .p2_2_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_2_2_ce0),
        .p2_2_2_q0(p2_2_2_q0),
        .p2_3_0_address0(grp_pointsOverlap_double_s_fu_238_p2_3_0_address0),
        .p2_3_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_3_0_ce0),
        .p2_3_0_q0(p2_3_0_q0),
        .p2_3_1_address0(grp_pointsOverlap_double_s_fu_238_p2_3_1_address0),
        .p2_3_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_3_1_ce0),
        .p2_3_1_q0(p2_3_1_q0),
        .p2_3_2_address0(grp_pointsOverlap_double_s_fu_238_p2_3_2_address0),
        .p2_3_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_3_2_ce0),
        .p2_3_2_q0(p2_3_2_q0),
        .p2_4_0_address0(grp_pointsOverlap_double_s_fu_238_p2_4_0_address0),
        .p2_4_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_4_0_ce0),
        .p2_4_0_q0(p2_4_0_q0),
        .p2_4_1_address0(grp_pointsOverlap_double_s_fu_238_p2_4_1_address0),
        .p2_4_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_4_1_ce0),
        .p2_4_1_q0(p2_4_1_q0),
        .p2_4_2_address0(grp_pointsOverlap_double_s_fu_238_p2_4_2_address0),
        .p2_4_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_4_2_ce0),
        .p2_4_2_q0(p2_4_2_q0),
        .p2_5_0_address0(grp_pointsOverlap_double_s_fu_238_p2_5_0_address0),
        .p2_5_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_5_0_ce0),
        .p2_5_0_q0(p2_5_0_q0),
        .p2_5_1_address0(grp_pointsOverlap_double_s_fu_238_p2_5_1_address0),
        .p2_5_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_5_1_ce0),
        .p2_5_1_q0(p2_5_1_q0),
        .p2_5_2_address0(grp_pointsOverlap_double_s_fu_238_p2_5_2_address0),
        .p2_5_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_5_2_ce0),
        .p2_5_2_q0(p2_5_2_q0),
        .p2_6_0_address0(grp_pointsOverlap_double_s_fu_238_p2_6_0_address0),
        .p2_6_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_6_0_ce0),
        .p2_6_0_q0(p2_6_0_q0),
        .p2_6_1_address0(grp_pointsOverlap_double_s_fu_238_p2_6_1_address0),
        .p2_6_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_6_1_ce0),
        .p2_6_1_q0(p2_6_1_q0),
        .p2_6_2_address0(grp_pointsOverlap_double_s_fu_238_p2_6_2_address0),
        .p2_6_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_6_2_ce0),
        .p2_6_2_q0(p2_6_2_q0),
        .p2_7_0_address0(grp_pointsOverlap_double_s_fu_238_p2_7_0_address0),
        .p2_7_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_7_0_ce0),
        .p2_7_0_q0(p2_7_0_q0),
        .p2_7_1_address0(grp_pointsOverlap_double_s_fu_238_p2_7_1_address0),
        .p2_7_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_7_1_ce0),
        .p2_7_1_q0(p2_7_1_q0),
        .p2_7_2_address0(grp_pointsOverlap_double_s_fu_238_p2_7_2_address0),
        .p2_7_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_7_2_ce0),
        .p2_7_2_q0(p2_7_2_q0),
        .p2_8_0_address0(grp_pointsOverlap_double_s_fu_238_p2_8_0_address0),
        .p2_8_0_ce0(grp_pointsOverlap_double_s_fu_238_p2_8_0_ce0),
        .p2_8_0_q0(p2_8_0_q0),
        .p2_8_1_address0(grp_pointsOverlap_double_s_fu_238_p2_8_1_address0),
        .p2_8_1_ce0(grp_pointsOverlap_double_s_fu_238_p2_8_1_ce0),
        .p2_8_1_q0(p2_8_1_q0),
        .p2_8_2_address0(grp_pointsOverlap_double_s_fu_238_p2_8_2_address0),
        .p2_8_2_ce0(grp_pointsOverlap_double_s_fu_238_p2_8_2_ce0),
        .p2_8_2_q0(p2_8_2_q0),
        .p2_offset(p2_offset),
        .p_read(cm_0_reg_711),
        .p_read1(cm_1_reg_716),
        .p_read2(cm_2_reg_721),
        .ap_return(grp_pointsOverlap_double_s_fu_238_ap_return)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage76),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_state77) & (ap_loop_exit_ready == 1'b1))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg <= 1'd0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state77) & ((icmp_ln184_reg_573 == 1'd1) | (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd0)))) begin
                ap_return_preg <= ap_phi_mux_merge_phi_fu_230_p4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_pointsOverlap_double_s_fu_238_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_NS_fsm_state19) & (1'b1 == ap_CS_fsm_state18) & (icmp_ln184_reg_573 == 1'd0))) begin
                grp_pointsOverlap_double_s_fu_238_ap_start_reg <= 1'b1;
            end else if ((grp_pointsOverlap_double_s_fu_238_ap_ready == 1'b1)) begin
                grp_pointsOverlap_double_s_fu_238_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            i_3_fu_128 <= 2'd0;
        end else if (((1'b1 == ap_CS_fsm_state77) & (icmp_ln184_reg_573 == 1'd0) & (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd1))) begin
            i_3_fu_128 <= select_ln184_2_fu_513_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            indvar_flatten_fu_132 <= 4'd0;
        end else if (((1'b1 == ap_CS_fsm_state77) & (icmp_ln184_reg_573 == 1'd0) & (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd1))) begin
            indvar_flatten_fu_132 <= add_ln184_3_reg_577;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            j_fu_124 <= 2'd0;
        end else if (((1'b1 == ap_CS_fsm_state77) & (icmp_ln184_reg_573 == 1'd0) & (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd1))) begin
            j_fu_124 <= add_ln185_fu_518_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state77) & (icmp_ln184_reg_573 == 1'd0) & (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd0))) begin
            merge_reg_226 <= 1'd0;
        end else if (((icmp_ln184_fu_378_p2 == 1'd1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            merge_reg_226 <= 1'd1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            add_ln179_reg_604 <= add_ln179_fu_447_p2;
            add_ln184_3_reg_577 <= add_ln184_3_fu_384_p2;
            add_ln184_reg_582 <= add_ln184_fu_393_p2;
            i_reg_568 <= ap_sig_allocacmp_i;
            icmp_ln184_reg_573 <= icmp_ln184_fu_378_p2;
            icmp_ln185_reg_587 <= icmp_ln185_fu_399_p2;
            select_ln184_1_reg_597 <= select_ln184_1_fu_435_p3;
            select_ln184_reg_592 <= select_ln184_fu_405_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            axes1_load_1_reg_641 <= axes1_q0;
            axes1_load_reg_635   <= axes1_q1;
            axes2_load_1_reg_663 <= axes2_q0;
            axes2_load_reg_657   <= axes2_q1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            axes1_load_2_reg_669 <= axes1_q0;
            axes2_load_2_reg_675 <= axes2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            cm_0_reg_711 <= grp_fu_469_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state18)) begin
            cm_1_reg_716 <= grp_fu_469_p_dout0;
            cm_2_reg_721 <= grp_fu_473_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            mul12_i_reg_696 <= grp_fu_497_p_dout0;
            mul17_i_reg_701 <= grp_fu_501_p_dout0;
            mul20_i_reg_706 <= grp_fu_505_p_dout0;
            mul9_i_reg_691  <= grp_fu_493_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            mul5_i_reg_686 <= grp_fu_497_p_dout0;
            mul_i_reg_681  <= grp_fu_493_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            sub_ln179_1_reg_620 <= sub_ln179_1_fu_478_p2;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state1_pp0_stage0_iter0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    assign ap_ST_fsm_state73_blk = 1'b0;

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state75_blk = 1'b0;

    assign ap_ST_fsm_state76_blk = 1'b0;

    assign ap_ST_fsm_state77_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state77) & ((icmp_ln184_reg_573 == 1'd1) | (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd0)))) begin
            ap_condition_exit_pp0_iter0_stage76 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage76 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state77) & (ap_loop_exit_ready == 1'b1))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state77) & (icmp_ln184_reg_573 == 1'd0) & (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd0))) begin
            ap_phi_mux_merge_phi_fu_230_p4 = 1'd0;
        end else begin
            ap_phi_mux_merge_phi_fu_230_p4 = merge_reg_226;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state77)) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state77) & ((icmp_ln184_reg_573 == 1'd1) | (grp_pointsOverlap_double_s_fu_238_ap_return == 1'd0)))) begin
            ap_return = ap_phi_mux_merge_phi_fu_230_p4;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_sig_allocacmp_i = 2'd0;
        end else begin
            ap_sig_allocacmp_i = i_3_fu_128;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_sig_allocacmp_indvar_flatten_load = 4'd0;
        end else begin
            ap_sig_allocacmp_indvar_flatten_load = indvar_flatten_fu_132;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_sig_allocacmp_j_load = 2'd0;
        end else begin
            ap_sig_allocacmp_j_load = j_fu_124;
        end
    end

    always @(*) begin
        if ((icmp_ln184_reg_573 == 1'd0)) begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                axes1_address0 = zext_ln184_fu_505_p1;
            end else if ((1'b1 == ap_CS_fsm_state2)) begin
                axes1_address0 = add_ln184_2_cast_fu_468_p1;
            end else begin
                axes1_address0 = 'bx;
            end
        end else begin
            axes1_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b1 == ap_CS_fsm_state3) & (icmp_ln184_reg_573 == 1'd0)) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln184_reg_573 == 1'd0)))) begin
            axes1_ce0 = 1'b1;
        end else begin
            axes1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            axes1_ce1 = 1'b1;
        end else begin
            axes1_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((icmp_ln184_reg_573 == 1'd0)) begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                axes2_address0 = zext_ln179_1_fu_509_p1;
            end else if ((1'b1 == ap_CS_fsm_state2)) begin
                axes2_address0 = zext_ln179_3_fu_500_p1;
            end else begin
                axes2_address0 = 'bx;
            end
        end else begin
            axes2_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b1 == ap_CS_fsm_state3) & (icmp_ln184_reg_573 == 1'd0)) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln184_reg_573 == 1'd0)))) begin
            axes2_ce0 = 1'b1;
        end else begin
            axes2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            axes2_ce1 = 1'b1;
        end else begin
            axes2_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_303_p0 = mul9_i_reg_691;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_303_p0 = mul_i_reg_681;
        end else begin
            grp_fu_303_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_303_p1 = mul12_i_reg_696;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_303_p1 = mul5_i_reg_686;
        end else begin
            grp_fu_303_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_311_p0 = axes1_load_1_reg_641;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_311_p0 = axes1_load_reg_635;
        end else begin
            grp_fu_311_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_311_p1 = axes2_load_2_reg_675;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_311_p1 = axes2_load_reg_657;
        end else begin
            grp_fu_311_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_315_p0 = axes1_load_2_reg_669;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_315_p0 = axes1_load_1_reg_641;
        end else begin
            grp_fu_315_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            grp_fu_315_p1 = axes2_load_reg_657;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_315_p1 = axes2_load_1_reg_663;
        end else begin
            grp_fu_315_p1 = 'bx;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln179_1_fu_483_p2 = (sub_ln179_1_fu_478_p2 + 7'd2);

    assign add_ln179_2_fu_494_p2 = (sub_ln179_1_fu_478_p2 + 7'd1);

    assign add_ln179_fu_447_p2 = ($signed(
        sub_ln179_cast_fu_327_p1
    ) + $signed(
        zext_ln179_fu_443_p1
    ));

    assign add_ln184_1_cast_fu_458_p1 = add_ln184_1_fu_453_p2;

    assign add_ln184_1_fu_453_p2 = (select_ln184_1_reg_597 + 6'd1);

    assign add_ln184_2_cast_fu_468_p1 = add_ln184_2_fu_463_p2;

    assign add_ln184_2_fu_463_p2 = (select_ln184_1_reg_597 + 6'd2);

    assign add_ln184_3_fu_384_p2 = (ap_sig_allocacmp_indvar_flatten_load + 4'd1);

    assign add_ln184_cast_fu_413_p1 = add_ln184_fu_393_p2;

    assign add_ln184_fu_393_p2 = (ap_sig_allocacmp_i + 2'd1);

    assign add_ln185_fu_518_p2 = (select_ln184_reg_592 + 2'd1);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

    assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];

    assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];

    assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state77 = ap_CS_fsm[32'd76];

    assign ap_NS_fsm_state19 = ap_NS_fsm[32'd18];

    always @(*) begin
        ap_block_state1_pp0_stage0_iter0 = (ap_start_int == 1'b0);
    end

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage76;

    assign axes1_address1 = add_ln184_1_cast_fu_458_p1;

    assign axes2_address1 = zext_ln179_2_fu_489_p1;

    assign empty_80_fu_360_p2 = ($signed(p_cast_fu_331_p1) + $signed(i_3_cast_fu_356_p1));

    assign empty_81_fu_366_p2 = empty_80_fu_360_p2 << 6'd2;

    assign empty_82_fu_372_p2 = (empty_81_fu_366_p2 - empty_80_fu_360_p2);

    assign empty_83_fu_417_p2 = ($signed(p_cast_fu_331_p1) + $signed(add_ln184_cast_fu_413_p1));

    assign empty_84_fu_423_p2 = empty_83_fu_417_p2 << 6'd2;

    assign empty_85_fu_429_p2 = (empty_84_fu_423_p2 - empty_83_fu_417_p2);

    assign grp_fu_469_p_ce = 1'b1;

    assign grp_fu_469_p_din0 = grp_fu_303_p0;

    assign grp_fu_469_p_din1 = grp_fu_303_p1;

    assign grp_fu_469_p_opcode = 2'd1;

    assign grp_fu_473_p_ce = 1'b1;

    assign grp_fu_473_p_din0 = mul17_i_reg_701;

    assign grp_fu_473_p_din1 = mul20_i_reg_706;

    assign grp_fu_473_p_opcode = 2'd1;

    assign grp_fu_493_p_ce = 1'b1;

    assign grp_fu_493_p_din0 = grp_fu_311_p0;

    assign grp_fu_493_p_din1 = grp_fu_311_p1;

    assign grp_fu_497_p_ce = 1'b1;

    assign grp_fu_497_p_din0 = grp_fu_315_p0;

    assign grp_fu_497_p_din1 = grp_fu_315_p1;

    assign grp_fu_501_p_ce = 1'b1;

    assign grp_fu_501_p_din0 = axes1_load_2_reg_669;

    assign grp_fu_501_p_din1 = axes2_load_1_reg_663;

    assign grp_fu_505_p_ce = 1'b1;

    assign grp_fu_505_p_din0 = axes1_load_reg_635;

    assign grp_fu_505_p_din1 = axes2_load_2_reg_675;

    assign grp_pointsOverlap_double_s_fu_238_ap_start = grp_pointsOverlap_double_s_fu_238_ap_start_reg;

    assign i_3_cast_fu_356_p1 = ap_sig_allocacmp_i;

    assign icmp_ln184_fu_378_p2 = ((ap_sig_allocacmp_indvar_flatten_load == 4'd9) ? 1'b1 : 1'b0);

    assign icmp_ln185_fu_399_p2 = ((ap_sig_allocacmp_j_load == 2'd3) ? 1'b1 : 1'b0);

    assign p1_address0 = grp_pointsOverlap_double_s_fu_238_p1_address0;

    assign p1_address1 = grp_pointsOverlap_double_s_fu_238_p1_address1;

    assign p1_ce0 = grp_pointsOverlap_double_s_fu_238_p1_ce0;

    assign p1_ce1 = grp_pointsOverlap_double_s_fu_238_p1_ce1;

    assign p2_0_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_0_0_address0;

    assign p2_0_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_0_0_ce0;

    assign p2_0_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_0_1_address0;

    assign p2_0_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_0_1_ce0;

    assign p2_0_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_0_2_address0;

    assign p2_0_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_0_2_ce0;

    assign p2_1_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_1_0_address0;

    assign p2_1_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_1_0_ce0;

    assign p2_1_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_1_1_address0;

    assign p2_1_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_1_1_ce0;

    assign p2_1_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_1_2_address0;

    assign p2_1_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_1_2_ce0;

    assign p2_2_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_2_0_address0;

    assign p2_2_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_2_0_ce0;

    assign p2_2_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_2_1_address0;

    assign p2_2_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_2_1_ce0;

    assign p2_2_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_2_2_address0;

    assign p2_2_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_2_2_ce0;

    assign p2_3_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_3_0_address0;

    assign p2_3_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_3_0_ce0;

    assign p2_3_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_3_1_address0;

    assign p2_3_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_3_1_ce0;

    assign p2_3_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_3_2_address0;

    assign p2_3_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_3_2_ce0;

    assign p2_4_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_4_0_address0;

    assign p2_4_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_4_0_ce0;

    assign p2_4_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_4_1_address0;

    assign p2_4_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_4_1_ce0;

    assign p2_4_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_4_2_address0;

    assign p2_4_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_4_2_ce0;

    assign p2_5_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_5_0_address0;

    assign p2_5_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_5_0_ce0;

    assign p2_5_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_5_1_address0;

    assign p2_5_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_5_1_ce0;

    assign p2_5_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_5_2_address0;

    assign p2_5_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_5_2_ce0;

    assign p2_6_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_6_0_address0;

    assign p2_6_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_6_0_ce0;

    assign p2_6_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_6_1_address0;

    assign p2_6_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_6_1_ce0;

    assign p2_6_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_6_2_address0;

    assign p2_6_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_6_2_ce0;

    assign p2_7_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_7_0_address0;

    assign p2_7_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_7_0_ce0;

    assign p2_7_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_7_1_address0;

    assign p2_7_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_7_1_ce0;

    assign p2_7_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_7_2_address0;

    assign p2_7_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_7_2_ce0;

    assign p2_8_0_address0 = grp_pointsOverlap_double_s_fu_238_p2_8_0_address0;

    assign p2_8_0_ce0 = grp_pointsOverlap_double_s_fu_238_p2_8_0_ce0;

    assign p2_8_1_address0 = grp_pointsOverlap_double_s_fu_238_p2_8_1_address0;

    assign p2_8_1_ce0 = grp_pointsOverlap_double_s_fu_238_p2_8_1_ce0;

    assign p2_8_2_address0 = grp_pointsOverlap_double_s_fu_238_p2_8_2_address0;

    assign p2_8_2_ce0 = grp_pointsOverlap_double_s_fu_238_p2_8_2_ce0;

    assign p_cast_fu_331_p1 = $signed(empty);

    assign select_ln184_1_fu_435_p3 = ((icmp_ln185_fu_399_p2[0:0] == 1'b1) ? empty_85_fu_429_p2 : empty_82_fu_372_p2);

    assign select_ln184_2_fu_513_p3 = ((icmp_ln185_reg_587[0:0] == 1'b1) ? add_ln184_reg_582 : i_reg_568);

    assign select_ln184_fu_405_p3 = ((icmp_ln185_fu_399_p2[0:0] == 1'b1) ? 2'd0 : ap_sig_allocacmp_j_load);

    assign shl_ln179_fu_473_p2 = add_ln179_reg_604 << 7'd2;

    assign sub_ln179_1_fu_478_p2 = (shl_ln179_fu_473_p2 - add_ln179_reg_604);

    assign sub_ln179_cast_fu_327_p1 = $signed(sub_ln179);

    assign zext_ln179_1_fu_509_p1 = sub_ln179_1_reg_620;

    assign zext_ln179_2_fu_489_p1 = add_ln179_1_fu_483_p2;

    assign zext_ln179_3_fu_500_p1 = add_ln179_2_fu_494_p2;

    assign zext_ln179_fu_443_p1 = select_ln184_fu_405_p3;

    assign zext_ln184_fu_505_p1 = select_ln184_1_reg_597;

endmodule  //main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_184_3_VITIS_LOOP_185_4
