/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_updateSensor (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    pf_address0,
    pf_ce0,
    pf_we0,
    pf_d0,
    pf_q0,
    pf_address1,
    pf_ce1,
    pf_q1,
    laserReading_address0,
    laserReading_ce0,
    laserReading_q0,
    laserReading_offset,
    grp_fu_401_p_din0,
    grp_fu_401_p_din1,
    grp_fu_401_p_opcode,
    grp_fu_401_p_dout0,
    grp_fu_401_p_ce,
    grp_fu_397_p_din0,
    grp_fu_397_p_din1,
    grp_fu_397_p_opcode,
    grp_fu_397_p_dout0,
    grp_fu_397_p_ce,
    grp_fu_405_p_din0,
    grp_fu_405_p_din1,
    grp_fu_405_p_dout0,
    grp_fu_405_p_ce,
    grp_fu_409_p_din0,
    grp_fu_409_p_din1,
    grp_fu_409_p_dout0,
    grp_fu_409_p_ce,
    grp_fu_394_p_din0,
    grp_fu_394_p_dout0,
    grp_fu_394_p_ce,
    grp_fu_413_p_din0,
    grp_fu_413_p_din1,
    grp_fu_413_p_opcode,
    grp_fu_413_p_dout0,
    grp_fu_413_p_ce,
    grp_fu_417_p_din0,
    grp_fu_417_p_din1,
    grp_fu_417_p_dout0,
    grp_fu_417_p_ce,
    grp_sin_or_cos_double_s_fu_421_p_din1,
    grp_sin_or_cos_double_s_fu_421_p_din2,
    grp_sin_or_cos_double_s_fu_421_p_dout0,
    grp_sin_or_cos_double_s_fu_421_p_start,
    grp_sin_or_cos_double_s_fu_421_p_ready,
    grp_sin_or_cos_double_s_fu_421_p_done,
    grp_sin_or_cos_double_s_fu_421_p_idle,
    grp_sin_or_cos_double_s_fu_432_p_din1,
    grp_sin_or_cos_double_s_fu_432_p_din2,
    grp_sin_or_cos_double_s_fu_432_p_dout0,
    grp_sin_or_cos_double_s_fu_432_p_start,
    grp_sin_or_cos_double_s_fu_432_p_ready,
    grp_sin_or_cos_double_s_fu_432_p_done,
    grp_sin_or_cos_double_s_fu_432_p_idle
);

    parameter ap_ST_fsm_state1 = 74'd1;
    parameter ap_ST_fsm_state2 = 74'd2;
    parameter ap_ST_fsm_state3 = 74'd4;
    parameter ap_ST_fsm_state4 = 74'd8;
    parameter ap_ST_fsm_state5 = 74'd16;
    parameter ap_ST_fsm_state6 = 74'd32;
    parameter ap_ST_fsm_state7 = 74'd64;
    parameter ap_ST_fsm_state8 = 74'd128;
    parameter ap_ST_fsm_state9 = 74'd256;
    parameter ap_ST_fsm_state10 = 74'd512;
    parameter ap_ST_fsm_state11 = 74'd1024;
    parameter ap_ST_fsm_state12 = 74'd2048;
    parameter ap_ST_fsm_state13 = 74'd4096;
    parameter ap_ST_fsm_state14 = 74'd8192;
    parameter ap_ST_fsm_state15 = 74'd16384;
    parameter ap_ST_fsm_state16 = 74'd32768;
    parameter ap_ST_fsm_state17 = 74'd65536;
    parameter ap_ST_fsm_state18 = 74'd131072;
    parameter ap_ST_fsm_state19 = 74'd262144;
    parameter ap_ST_fsm_state20 = 74'd524288;
    parameter ap_ST_fsm_state21 = 74'd1048576;
    parameter ap_ST_fsm_state22 = 74'd2097152;
    parameter ap_ST_fsm_state23 = 74'd4194304;
    parameter ap_ST_fsm_state24 = 74'd8388608;
    parameter ap_ST_fsm_state25 = 74'd16777216;
    parameter ap_ST_fsm_state26 = 74'd33554432;
    parameter ap_ST_fsm_state27 = 74'd67108864;
    parameter ap_ST_fsm_state28 = 74'd134217728;
    parameter ap_ST_fsm_state29 = 74'd268435456;
    parameter ap_ST_fsm_state30 = 74'd536870912;
    parameter ap_ST_fsm_state31 = 74'd1073741824;
    parameter ap_ST_fsm_state32 = 74'd2147483648;
    parameter ap_ST_fsm_state33 = 74'd4294967296;
    parameter ap_ST_fsm_state34 = 74'd8589934592;
    parameter ap_ST_fsm_state35 = 74'd17179869184;
    parameter ap_ST_fsm_state36 = 74'd34359738368;
    parameter ap_ST_fsm_state37 = 74'd68719476736;
    parameter ap_ST_fsm_state38 = 74'd137438953472;
    parameter ap_ST_fsm_state39 = 74'd274877906944;
    parameter ap_ST_fsm_state40 = 74'd549755813888;
    parameter ap_ST_fsm_state41 = 74'd1099511627776;
    parameter ap_ST_fsm_state42 = 74'd2199023255552;
    parameter ap_ST_fsm_state43 = 74'd4398046511104;
    parameter ap_ST_fsm_state44 = 74'd8796093022208;
    parameter ap_ST_fsm_state45 = 74'd17592186044416;
    parameter ap_ST_fsm_state46 = 74'd35184372088832;
    parameter ap_ST_fsm_state47 = 74'd70368744177664;
    parameter ap_ST_fsm_state48 = 74'd140737488355328;
    parameter ap_ST_fsm_state49 = 74'd281474976710656;
    parameter ap_ST_fsm_state50 = 74'd562949953421312;
    parameter ap_ST_fsm_state51 = 74'd1125899906842624;
    parameter ap_ST_fsm_state52 = 74'd2251799813685248;
    parameter ap_ST_fsm_state53 = 74'd4503599627370496;
    parameter ap_ST_fsm_state54 = 74'd9007199254740992;
    parameter ap_ST_fsm_state55 = 74'd18014398509481984;
    parameter ap_ST_fsm_state56 = 74'd36028797018963968;
    parameter ap_ST_fsm_state57 = 74'd72057594037927936;
    parameter ap_ST_fsm_state58 = 74'd144115188075855872;
    parameter ap_ST_fsm_state59 = 74'd288230376151711744;
    parameter ap_ST_fsm_state60 = 74'd576460752303423488;
    parameter ap_ST_fsm_state61 = 74'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 74'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 74'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 74'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 74'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 74'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 74'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 74'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 74'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 74'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 74'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 74'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 74'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 74'd9444732965739290427392;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [16:0] pf_address0;
    output pf_ce0;
    output [31:0] pf_we0;
    output [255:0] pf_d0;
    input [255:0] pf_q0;
    output [16:0] pf_address1;
    output pf_ce1;
    input [255:0] pf_q1;
    output [17:0] laserReading_address0;
    output laserReading_ce0;
    input [31:0] laserReading_q0;
    input [9:0] laserReading_offset;
    output [63:0] grp_fu_401_p_din0;
    output [63:0] grp_fu_401_p_din1;
    output [1:0] grp_fu_401_p_opcode;
    input [63:0] grp_fu_401_p_dout0;
    output grp_fu_401_p_ce;
    output [63:0] grp_fu_397_p_din0;
    output [63:0] grp_fu_397_p_din1;
    output [0:0] grp_fu_397_p_opcode;
    input [63:0] grp_fu_397_p_dout0;
    output grp_fu_397_p_ce;
    output [63:0] grp_fu_405_p_din0;
    output [63:0] grp_fu_405_p_din1;
    input [63:0] grp_fu_405_p_dout0;
    output grp_fu_405_p_ce;
    output [63:0] grp_fu_409_p_din0;
    output [63:0] grp_fu_409_p_din1;
    input [63:0] grp_fu_409_p_dout0;
    output grp_fu_409_p_ce;
    output [31:0] grp_fu_394_p_din0;
    input [63:0] grp_fu_394_p_dout0;
    output grp_fu_394_p_ce;
    output [63:0] grp_fu_413_p_din0;
    output [63:0] grp_fu_413_p_din1;
    output [4:0] grp_fu_413_p_opcode;
    input [0:0] grp_fu_413_p_dout0;
    output grp_fu_413_p_ce;
    output [63:0] grp_fu_417_p_din0;
    output [63:0] grp_fu_417_p_din1;
    input [63:0] grp_fu_417_p_dout0;
    output grp_fu_417_p_ce;
    output [63:0] grp_sin_or_cos_double_s_fu_421_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_421_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_421_p_dout0;
    output grp_sin_or_cos_double_s_fu_421_p_start;
    input grp_sin_or_cos_double_s_fu_421_p_ready;
    input grp_sin_or_cos_double_s_fu_421_p_done;
    input grp_sin_or_cos_double_s_fu_421_p_idle;
    output [63:0] grp_sin_or_cos_double_s_fu_432_p_din1;
    output [0:0] grp_sin_or_cos_double_s_fu_432_p_din2;
    input [63:0] grp_sin_or_cos_double_s_fu_432_p_dout0;
    output grp_sin_or_cos_double_s_fu_432_p_start;
    input grp_sin_or_cos_double_s_fu_432_p_ready;
    input grp_sin_or_cos_double_s_fu_432_p_done;
    input grp_sin_or_cos_double_s_fu_432_p_idle;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[16:0] pf_address0;
    reg pf_ce0;
    reg[31:0] pf_we0;
    reg[16:0] pf_address1;
    reg pf_ce1;

    (* fsm_encoding = "none" *) reg   [73:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire   [17:0] mul_ln177_fu_253_p2;
    reg   [17:0] mul_ln177_reg_444;
    wire   [8:0] add_ln162_fu_273_p2;
    reg   [8:0] add_ln162_reg_467;
    wire    ap_CS_fsm_state2;
    reg   [16:0] pf_addr_3_reg_472;
    wire   [63:0] x_fu_288_p1;
    reg   [63:0] x_reg_478;
    wire    ap_CS_fsm_state3;
    wire   [63:0] y_fu_292_p1;
    reg   [63:0] y_reg_483;
    wire   [63:0] theta_fu_296_p1;
    reg   [63:0] theta_reg_488;
    reg   [17:0] trunc_ln3_reg_493;
    wire  signed [32:0] sext_ln168_fu_320_p1;
    reg  signed [32:0] sext_ln168_reg_498;
    wire    ap_CS_fsm_state4;
    wire   [32:0] add_ln168_fu_335_p2;
    reg   [32:0] add_ln168_reg_511;
    wire   [63:0] grp_fu_226_p1;
    reg   [63:0] conv_reg_516;
    wire    ap_CS_fsm_state9;
    wire   [254:0] empty_fu_349_p1;
    reg   [254:0] empty_reg_521;
    wire    ap_CS_fsm_state12;
    reg   [63:0] p_cast2_reg_526;
    wire   [63:0] trunc_ln205_fu_363_p1;
    reg   [63:0] trunc_ln205_reg_531;
    reg   [51:0] trunc_ln188_2_reg_536;
    wire   [63:0] empty_64_fu_377_p1;
    reg   [63:0] empty_64_reg_541;
    wire    ap_CS_fsm_state13;
    wire   [63:0] grp_fu_221_p2;
    reg   [63:0] pRand_reg_547;
    wire    ap_CS_fsm_state71;
    wire   [63:0] empty_65_fu_381_p1;
    reg   [63:0] empty_65_reg_552;
    wire   [63:0] grp_fu_229_p4;
    reg   [63:0] p_cast4_reg_557;
    wire   [63:0] grp_fu_239_p4;
    reg   [63:0] p_cast6_reg_562;
    reg   [63:0] p_cast7_reg_567;
    wire   [63:0] empty_66_fu_395_p1;
    reg   [63:0] empty_66_reg_572;
    wire    ap_CS_fsm_state72;
    wire   [63:0] empty_67_fu_399_p1;
    reg   [63:0] empty_67_reg_577;
    wire   [63:0] empty_68_fu_403_p1;
    reg   [63:0] empty_68_reg_582;
    wire   [63:0] empty_69_fu_407_p1;
    reg   [63:0] empty_69_reg_587;
    wire   [63:0] bitcast_ln205_fu_411_p1;
    reg   [63:0] bitcast_ln205_reg_592;
    reg   [7:0] zStar_address0;
    reg    zStar_ce0;
    reg    zStar_we0;
    wire   [63:0] zStar_q0;
    wire    grp_rayCast_fu_179_ap_start;
    wire    grp_rayCast_fu_179_ap_done;
    wire    grp_rayCast_fu_179_ap_idle;
    wire    grp_rayCast_fu_179_ap_ready;
    wire   [16:0] grp_rayCast_fu_179_pf_address0;
    wire    grp_rayCast_fu_179_pf_ce0;
    wire   [63:0] grp_rayCast_fu_179_ap_return;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_597_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_597_p_din1;
    wire   [1:0] grp_rayCast_fu_179_grp_fu_597_p_opcode;
    wire    grp_rayCast_fu_179_grp_fu_597_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_601_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_601_p_din1;
    wire   [0:0] grp_rayCast_fu_179_grp_fu_601_p_opcode;
    wire    grp_rayCast_fu_179_grp_fu_601_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_605_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_605_p_din1;
    wire    grp_rayCast_fu_179_grp_fu_605_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_609_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_609_p_din1;
    wire    grp_rayCast_fu_179_grp_fu_609_p_ce;
    wire   [31:0] grp_rayCast_fu_179_grp_fu_613_p_din0;
    wire    grp_rayCast_fu_179_grp_fu_613_p_ce;
    wire   [31:0] grp_rayCast_fu_179_grp_fu_616_p_din0;
    wire   [31:0] grp_rayCast_fu_179_grp_fu_616_p_din1;
    wire   [4:0] grp_rayCast_fu_179_grp_fu_616_p_opcode;
    wire    grp_rayCast_fu_179_grp_fu_616_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_221_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_221_p_din1;
    wire    grp_rayCast_fu_179_grp_fu_221_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_620_p_din0;
    wire   [63:0] grp_rayCast_fu_179_grp_fu_620_p_din1;
    wire   [4:0] grp_rayCast_fu_179_grp_fu_620_p_opcode;
    wire    grp_rayCast_fu_179_grp_fu_620_p_ce;
    wire   [63:0] grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din1;
    wire  signed [0:0] grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din2;
    wire    grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_start;
    wire   [63:0] grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din1;
    wire   [0:0] grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din2;
    wire    grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_start;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_done;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_idle;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_ready;
    wire   [17:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_address0;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_ce0;
    wire   [7:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_address0;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_ce0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_probability_out;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_probability_out_ap_vld;
    wire   [31:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_din0;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_ce;
    wire   [31:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din0;
    wire   [31:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din1;
    wire   [4:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_opcode;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din1;
    wire   [1:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_opcode;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din1;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din1;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din1;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din1;
    wire   [4:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_opcode;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_ce;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din0;
    wire   [63:0] grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din1;
    wire    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_ce;
    reg    grp_sin_or_cos_double_s_fu_624_ap_start;
    reg    grp_sin_or_cos_double_s_fu_635_ap_start;
    reg   [32:0] d_reg_167;
    wire    ap_CS_fsm_state11;
    reg    grp_rayCast_fu_179_ap_start_reg;
    wire    ap_CS_fsm_state10;
    reg    grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg;
    wire    ap_CS_fsm_state73;
    wire   [63:0] zext_ln162_fu_279_p1;
    wire   [0:0] icmp_ln162_fu_267_p2;
    wire   [63:0] zext_ln168_fu_344_p1;
    reg   [8:0] i_fu_96;
    wire   [0:0] icmp_ln168_fu_324_p2;
    wire    ap_CS_fsm_state74;
    wire    ap_CS_fsm_state70;
    reg   [63:0] grp_fu_221_p0;
    reg   [63:0] grp_fu_221_p1;
    wire   [31:0] grp_fu_226_p0;
    wire   [9:0] mul_ln177_fu_253_p0;
    wire   [8:0] mul_ln177_fu_253_p1;
    wire   [63:0] trunc_ln163_fu_284_p1;
    wire   [31:0] p_cast_fu_300_p4;
    wire   [63:0] bitcast_ln181_fu_418_p1;
    reg    grp_fu_221_ce;
    reg   [63:0] grp_fu_597_p0;
    reg   [63:0] grp_fu_597_p1;
    reg   [1:0] grp_fu_597_opcode;
    reg    grp_fu_597_ce;
    reg    grp_fu_601_ce;
    reg   [63:0] grp_fu_605_p0;
    reg   [63:0] grp_fu_605_p1;
    reg    grp_fu_605_ce;
    reg   [63:0] grp_fu_609_p0;
    reg   [63:0] grp_fu_609_p1;
    reg    grp_fu_609_ce;
    reg   [31:0] grp_fu_613_p0;
    reg    grp_fu_613_ce;
    wire   [0:0] grp_fu_616_p2;
    reg   [31:0] grp_fu_616_p0;
    reg   [31:0] grp_fu_616_p1;
    reg    grp_fu_616_ce;
    reg   [4:0] grp_fu_616_opcode;
    reg   [63:0] grp_fu_620_p0;
    reg   [63:0] grp_fu_620_p1;
    reg    grp_fu_620_ce;
    reg   [4:0] grp_fu_620_opcode;
    reg    grp_fu_646_ce;
    reg   [73:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    reg    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_ST_fsm_state62_blk;
    wire    ap_ST_fsm_state63_blk;
    wire    ap_ST_fsm_state64_blk;
    wire    ap_ST_fsm_state65_blk;
    wire    ap_ST_fsm_state66_blk;
    wire    ap_ST_fsm_state67_blk;
    wire    ap_ST_fsm_state68_blk;
    wire    ap_ST_fsm_state69_blk;
    wire    ap_ST_fsm_state70_blk;
    wire    ap_ST_fsm_state71_blk;
    wire    ap_ST_fsm_state72_blk;
    reg    ap_ST_fsm_state73_blk;
    wire    ap_ST_fsm_state74_blk;
    wire   [17:0] mul_ln177_fu_253_p00;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 74'd1;
        #0 grp_rayCast_fu_179_ap_start_reg = 1'b0;
        #0 grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg = 1'b0;
        #0 i_fu_96 = 9'd0;
    end

    main_updateSensor_zStar_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(180),
        .AddressWidth(8)
    ) zStar_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(zStar_address0),
        .ce0(zStar_ce0),
        .we0(zStar_we0),
        .d0(grp_rayCast_fu_179_ap_return),
        .q0(zStar_q0)
    );

    main_rayCast grp_rayCast_fu_179 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_rayCast_fu_179_ap_start),
        .ap_done(grp_rayCast_fu_179_ap_done),
        .ap_idle(grp_rayCast_fu_179_ap_idle),
        .ap_ready(grp_rayCast_fu_179_ap_ready),
        .pf_address0(grp_rayCast_fu_179_pf_address0),
        .pf_ce0(grp_rayCast_fu_179_pf_ce0),
        .pf_q0(pf_q0),
        .x(x_reg_478),
        .y(y_reg_483),
        .theta(theta_reg_488),
        .degree(conv_reg_516),
        .ap_return(grp_rayCast_fu_179_ap_return),
        .grp_fu_597_p_din0(grp_rayCast_fu_179_grp_fu_597_p_din0),
        .grp_fu_597_p_din1(grp_rayCast_fu_179_grp_fu_597_p_din1),
        .grp_fu_597_p_opcode(grp_rayCast_fu_179_grp_fu_597_p_opcode),
        .grp_fu_597_p_dout0(grp_fu_401_p_dout0),
        .grp_fu_597_p_ce(grp_rayCast_fu_179_grp_fu_597_p_ce),
        .grp_fu_601_p_din0(grp_rayCast_fu_179_grp_fu_601_p_din0),
        .grp_fu_601_p_din1(grp_rayCast_fu_179_grp_fu_601_p_din1),
        .grp_fu_601_p_opcode(grp_rayCast_fu_179_grp_fu_601_p_opcode),
        .grp_fu_601_p_dout0(grp_fu_397_p_dout0),
        .grp_fu_601_p_ce(grp_rayCast_fu_179_grp_fu_601_p_ce),
        .grp_fu_605_p_din0(grp_rayCast_fu_179_grp_fu_605_p_din0),
        .grp_fu_605_p_din1(grp_rayCast_fu_179_grp_fu_605_p_din1),
        .grp_fu_605_p_dout0(grp_fu_405_p_dout0),
        .grp_fu_605_p_ce(grp_rayCast_fu_179_grp_fu_605_p_ce),
        .grp_fu_609_p_din0(grp_rayCast_fu_179_grp_fu_609_p_din0),
        .grp_fu_609_p_din1(grp_rayCast_fu_179_grp_fu_609_p_din1),
        .grp_fu_609_p_dout0(grp_fu_409_p_dout0),
        .grp_fu_609_p_ce(grp_rayCast_fu_179_grp_fu_609_p_ce),
        .grp_fu_613_p_din0(grp_rayCast_fu_179_grp_fu_613_p_din0),
        .grp_fu_613_p_dout0(grp_fu_394_p_dout0),
        .grp_fu_613_p_ce(grp_rayCast_fu_179_grp_fu_613_p_ce),
        .grp_fu_616_p_din0(grp_rayCast_fu_179_grp_fu_616_p_din0),
        .grp_fu_616_p_din1(grp_rayCast_fu_179_grp_fu_616_p_din1),
        .grp_fu_616_p_opcode(grp_rayCast_fu_179_grp_fu_616_p_opcode),
        .grp_fu_616_p_dout0(grp_fu_616_p2),
        .grp_fu_616_p_ce(grp_rayCast_fu_179_grp_fu_616_p_ce),
        .grp_fu_221_p_din0(grp_rayCast_fu_179_grp_fu_221_p_din0),
        .grp_fu_221_p_din1(grp_rayCast_fu_179_grp_fu_221_p_din1),
        .grp_fu_221_p_dout0(grp_fu_221_p2),
        .grp_fu_221_p_ce(grp_rayCast_fu_179_grp_fu_221_p_ce),
        .grp_fu_620_p_din0(grp_rayCast_fu_179_grp_fu_620_p_din0),
        .grp_fu_620_p_din1(grp_rayCast_fu_179_grp_fu_620_p_din1),
        .grp_fu_620_p_opcode(grp_rayCast_fu_179_grp_fu_620_p_opcode),
        .grp_fu_620_p_dout0(grp_fu_413_p_dout0),
        .grp_fu_620_p_ce(grp_rayCast_fu_179_grp_fu_620_p_ce),
        .grp_sin_or_cos_double_s_fu_624_p_din1(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din1),
        .grp_sin_or_cos_double_s_fu_624_p_din2(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din2),
        .grp_sin_or_cos_double_s_fu_624_p_dout0(grp_sin_or_cos_double_s_fu_421_p_dout0),
        .grp_sin_or_cos_double_s_fu_624_p_start(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_start),
        .grp_sin_or_cos_double_s_fu_624_p_ready(grp_sin_or_cos_double_s_fu_421_p_ready),
        .grp_sin_or_cos_double_s_fu_624_p_done(grp_sin_or_cos_double_s_fu_421_p_done),
        .grp_sin_or_cos_double_s_fu_624_p_idle(grp_sin_or_cos_double_s_fu_421_p_idle),
        .grp_sin_or_cos_double_s_fu_635_p_din1(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din1),
        .grp_sin_or_cos_double_s_fu_635_p_din2(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din2),
        .grp_sin_or_cos_double_s_fu_635_p_dout0(grp_sin_or_cos_double_s_fu_432_p_dout0),
        .grp_sin_or_cos_double_s_fu_635_p_start(grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_start),
        .grp_sin_or_cos_double_s_fu_635_p_ready(grp_sin_or_cos_double_s_fu_432_p_ready),
        .grp_sin_or_cos_double_s_fu_635_p_done(grp_sin_or_cos_double_s_fu_432_p_done),
        .grp_sin_or_cos_double_s_fu_635_p_idle(grp_sin_or_cos_double_s_fu_432_p_idle)
    );

    main_updateSensor_Pipeline_VITIS_LOOP_173_3 grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start),
        .ap_done(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_done),
        .ap_idle(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_idle),
        .ap_ready(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_ready),
        .empty_10(empty_66_reg_572),
        .empty_11(empty_67_reg_577),
        .empty_12(empty_68_reg_582),
        .empty_13(empty_69_reg_587),
        .empty(empty_64_reg_541),
        .trunc_ln3(trunc_ln3_reg_493),
        .mul_ln177(mul_ln177_reg_444),
        .laserReading_address0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_address0),
        .laserReading_ce0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_ce0),
        .laserReading_q0(laserReading_q0),
        .zStar_address0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_address0),
        .zStar_ce0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_ce0),
        .zStar_q0(zStar_q0),
        .pf_load_2(empty_reg_521),
        .trunc_ln188_2(trunc_ln188_2_reg_536),
        .pRand(pRand_reg_547),
        .bitcast_ln205(bitcast_ln205_reg_592),
        .probability_out(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_probability_out),
        .probability_out_ap_vld(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_probability_out_ap_vld),
        .grp_fu_613_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_din0),
        .grp_fu_613_p_dout0(grp_fu_394_p_dout0),
        .grp_fu_613_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_ce),
        .grp_fu_616_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din0),
        .grp_fu_616_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din1),
        .grp_fu_616_p_opcode(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_opcode),
        .grp_fu_616_p_dout0(grp_fu_616_p2),
        .grp_fu_616_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_ce),
        .grp_fu_597_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din0),
        .grp_fu_597_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din1),
        .grp_fu_597_p_opcode(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_opcode),
        .grp_fu_597_p_dout0(grp_fu_401_p_dout0),
        .grp_fu_597_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_ce),
        .grp_fu_605_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din0),
        .grp_fu_605_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din1),
        .grp_fu_605_p_dout0(grp_fu_405_p_dout0),
        .grp_fu_605_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_ce),
        .grp_fu_609_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din0),
        .grp_fu_609_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din1),
        .grp_fu_609_p_dout0(grp_fu_409_p_dout0),
        .grp_fu_609_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_ce),
        .grp_fu_221_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din0),
        .grp_fu_221_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din1),
        .grp_fu_221_p_dout0(grp_fu_221_p2),
        .grp_fu_221_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_ce),
        .grp_fu_620_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din0),
        .grp_fu_620_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din1),
        .grp_fu_620_p_opcode(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_opcode),
        .grp_fu_620_p_dout0(grp_fu_413_p_dout0),
        .grp_fu_620_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_ce),
        .grp_fu_646_p_din0(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din0),
        .grp_fu_646_p_din1(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din1),
        .grp_fu_646_p_dout0(grp_fu_417_p_dout0),
        .grp_fu_646_p_ce(grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_ce)
    );

    main_ddiv_64ns_64ns_64_59_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(59),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) ddiv_64ns_64ns_64_59_no_dsp_1_U194 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_221_p0),
        .din1(grp_fu_221_p1),
        .ce(grp_fu_221_ce),
        .dout(grp_fu_221_p2)
    );

    main_sitodp_32ns_64_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) sitodp_32ns_64_6_no_dsp_1_U195 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_226_p0),
        .ce(1'b1),
        .dout(grp_fu_226_p1)
    );

    main_mul_10ns_9ns_18_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(10),
        .din1_WIDTH(9),
        .dout_WIDTH(18)
    ) mul_10ns_9ns_18_1_1_U196 (
        .din0(mul_ln177_fu_253_p0),
        .din1(mul_ln177_fu_253_p1),
        .dout(mul_ln177_fu_253_p2)
    );

    main_fcmp_32ns_32ns_1_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(1)
    ) fcmp_32ns_32ns_1_2_no_dsp_1_U202 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_616_p0),
        .din1(grp_fu_616_p1),
        .ce(grp_fu_616_ce),
        .opcode(grp_fu_616_opcode),
        .dout(grp_fu_616_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_rayCast_fu_179_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state10)) begin
                grp_rayCast_fu_179_ap_start_reg <= 1'b1;
            end else if ((grp_rayCast_fu_179_ap_ready == 1'b1)) begin
                grp_rayCast_fu_179_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state72)) begin
                grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg <= 1'b1;
            end else if ((grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_ready == 1'b1)) begin
                grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            d_reg_167 <= 33'd0;
        end else if (((grp_rayCast_fu_179_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
            d_reg_167 <= add_ln168_reg_511;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            i_fu_96 <= 9'd0;
        end else if (((icmp_ln168_fu_324_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4))) begin
            i_fu_96 <= add_ln162_reg_467;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            add_ln162_reg_467 <= add_ln162_fu_273_p2;
            pf_addr_3_reg_472[8 : 0] <= zext_ln162_fu_279_p1[8 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            add_ln168_reg_511 <= add_ln168_fu_335_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state72)) begin
            bitcast_ln205_reg_592 <= bitcast_ln205_fu_411_p1;
            empty_66_reg_572 <= empty_66_fu_395_p1;
            empty_67_reg_577 <= empty_67_fu_399_p1;
            empty_68_reg_582 <= empty_68_fu_403_p1;
            empty_69_reg_587 <= empty_69_fu_407_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            conv_reg_516 <= grp_fu_226_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state13)) begin
            empty_64_reg_541 <= empty_64_fu_377_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state71)) begin
            empty_65_reg_552 <= empty_65_fu_381_p1;
            pRand_reg_547 <= grp_fu_221_p2;
            p_cast4_reg_557 <= {{pf_q1[127:64]}};
            p_cast6_reg_562 <= {{pf_q1[191:128]}};
            p_cast7_reg_567 <= {{pf_q1[255:192]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            empty_reg_521 <= empty_fu_349_p1;
            p_cast2_reg_526 <= {{pf_q0[255:192]}};
            trunc_ln188_2_reg_536 <= {{pf_q0[243:192]}};
            trunc_ln205_reg_531 <= trunc_ln205_fu_363_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            mul_ln177_reg_444 <= mul_ln177_fu_253_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            sext_ln168_reg_498 <= sext_ln168_fu_320_p1;
            theta_reg_488 <= theta_fu_296_p1;
            trunc_ln3_reg_493 <= {{pf_q0[145:128]}};
            x_reg_478 <= x_fu_288_p1;
            y_reg_483 <= y_fu_292_p1;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    always @(*) begin
        if ((grp_rayCast_fu_179_ap_done == 1'b0)) begin
            ap_ST_fsm_state11_blk = 1'b1;
        end else begin
            ap_ST_fsm_state11_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    always @(*) begin
        if ((grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_done == 1'b0)) begin
            ap_ST_fsm_state73_blk = 1'b1;
        end else begin
            ap_ST_fsm_state73_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if ((((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln162_fu_267_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln162_fu_267_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_221_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_221_ce = grp_rayCast_fu_179_grp_fu_221_p_ce;
        end else begin
            grp_fu_221_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_221_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_221_p0 = grp_rayCast_fu_179_grp_fu_221_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            grp_fu_221_p0 = 64'd4607182418800017408;
        end else begin
            grp_fu_221_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_221_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_221_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_221_p1 = grp_rayCast_fu_179_grp_fu_221_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            grp_fu_221_p1 = empty_64_fu_377_p1;
        end else begin
            grp_fu_221_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_597_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_597_ce = grp_rayCast_fu_179_grp_fu_597_p_ce;
        end else begin
            grp_fu_597_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_597_opcode = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_597_opcode = grp_rayCast_fu_179_grp_fu_597_p_opcode;
        end else begin
            grp_fu_597_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_597_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_597_p0 = grp_rayCast_fu_179_grp_fu_597_p_din0;
        end else begin
            grp_fu_597_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_597_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_597_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_597_p1 = grp_rayCast_fu_179_grp_fu_597_p_din1;
        end else begin
            grp_fu_597_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_601_ce = grp_rayCast_fu_179_grp_fu_601_p_ce;
        end else begin
            grp_fu_601_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_605_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_605_ce = grp_rayCast_fu_179_grp_fu_605_p_ce;
        end else begin
            grp_fu_605_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_605_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_605_p0 = grp_rayCast_fu_179_grp_fu_605_p_din0;
        end else begin
            grp_fu_605_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_605_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_605_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_605_p1 = grp_rayCast_fu_179_grp_fu_605_p_din1;
        end else begin
            grp_fu_605_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_609_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_609_ce = grp_rayCast_fu_179_grp_fu_609_p_ce;
        end else begin
            grp_fu_609_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_609_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_609_p0 = grp_rayCast_fu_179_grp_fu_609_p_din0;
        end else begin
            grp_fu_609_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_609_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_609_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_609_p1 = grp_rayCast_fu_179_grp_fu_609_p_din1;
        end else begin
            grp_fu_609_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_613_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_613_ce = grp_rayCast_fu_179_grp_fu_613_p_ce;
        end else begin
            grp_fu_613_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_613_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_613_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_613_p0 = grp_rayCast_fu_179_grp_fu_613_p_din0;
        end else begin
            grp_fu_613_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_616_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_616_ce = grp_rayCast_fu_179_grp_fu_616_p_ce;
        end else begin
            grp_fu_616_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_616_opcode = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_616_opcode = grp_rayCast_fu_179_grp_fu_616_p_opcode;
        end else begin
            grp_fu_616_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_616_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_616_p0 = grp_rayCast_fu_179_grp_fu_616_p_din0;
        end else begin
            grp_fu_616_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_616_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_616_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_616_p1 = grp_rayCast_fu_179_grp_fu_616_p_din1;
        end else begin
            grp_fu_616_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_620_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_620_ce = grp_rayCast_fu_179_grp_fu_620_p_ce;
        end else begin
            grp_fu_620_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_620_opcode = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_620_opcode = grp_rayCast_fu_179_grp_fu_620_p_opcode;
        end else begin
            grp_fu_620_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_620_p0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_620_p0 = grp_rayCast_fu_179_grp_fu_620_p_din0;
        end else begin
            grp_fu_620_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_620_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_620_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_620_p1 = grp_rayCast_fu_179_grp_fu_620_p_din1;
        end else begin
            grp_fu_620_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            grp_fu_646_ce = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_ce;
        end else begin
            grp_fu_646_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_sin_or_cos_double_s_fu_624_ap_start = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_start;
        end else begin
            grp_sin_or_cos_double_s_fu_624_ap_start = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_sin_or_cos_double_s_fu_635_ap_start = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_start;
        end else begin
            grp_sin_or_cos_double_s_fu_635_ap_start = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state74)) begin
            pf_address0 = pf_addr_3_reg_472;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            pf_address0 = 64'd80502;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            pf_address0 = 64'd80503;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            pf_address0 = grp_rayCast_fu_179_pf_address0;
        end else begin
            pf_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state70)) begin
            pf_address1 = 64'd80501;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            pf_address1 = zext_ln162_fu_279_p1;
        end else begin
            pf_address1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state2))) begin
            pf_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            pf_ce0 = grp_rayCast_fu_179_pf_ce0;
        end else begin
            pf_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state70) | (1'b1 == ap_CS_fsm_state2))) begin
            pf_ce1 = 1'b1;
        end else begin
            pf_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state74)) begin
            pf_we0 = 32'd4278190080;
        end else begin
            pf_we0 = 32'd0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            zStar_address0 = zext_ln168_fu_344_p1;
        end else if ((1'b1 == ap_CS_fsm_state73)) begin
            zStar_address0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_address0;
        end else begin
            zStar_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((grp_rayCast_fu_179_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
            zStar_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state73)) begin
            zStar_ce0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_zStar_ce0;
        end else begin
            zStar_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((grp_rayCast_fu_179_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
            zStar_we0 = 1'b1;
        end else begin
            zStar_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                if (((icmp_ln162_fu_267_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                if (((icmp_ln168_fu_324_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state4))) begin
                    ap_NS_fsm = ap_ST_fsm_state12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                if (((grp_rayCast_fu_179_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state11;
                end
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                if (((grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state73))) begin
                    ap_NS_fsm = ap_ST_fsm_state74;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state73;
                end
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln162_fu_273_p2 = (i_fu_96 + 9'd1);

    assign add_ln168_fu_335_p2 = ($signed(sext_ln168_reg_498) + $signed(d_reg_167));

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];

    assign ap_CS_fsm_state71 = ap_CS_fsm[32'd70];

    assign ap_CS_fsm_state72 = ap_CS_fsm[32'd71];

    assign ap_CS_fsm_state73 = ap_CS_fsm[32'd72];

    assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign bitcast_ln181_fu_418_p1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_probability_out;

    assign bitcast_ln205_fu_411_p1 = trunc_ln205_reg_531;

    assign empty_64_fu_377_p1 = p_cast2_reg_526;

    assign empty_65_fu_381_p1 = pf_q1[63:0];

    assign empty_66_fu_395_p1 = empty_65_reg_552;

    assign empty_67_fu_399_p1 = p_cast4_reg_557;

    assign empty_68_fu_403_p1 = p_cast6_reg_562;

    assign empty_69_fu_407_p1 = p_cast7_reg_567;

    assign empty_fu_349_p1 = pf_q0[254:0];

    assign grp_fu_226_p0 = d_reg_167[31:0];

    assign grp_fu_229_p4 = {{pf_q1[127:64]}};

    assign grp_fu_239_p4 = {{pf_q1[191:128]}};

    assign grp_fu_394_p_ce = grp_fu_613_ce;

    assign grp_fu_394_p_din0 = grp_fu_613_p0;

    assign grp_fu_397_p_ce = grp_fu_601_ce;

    assign grp_fu_397_p_din0 = grp_rayCast_fu_179_grp_fu_601_p_din0;

    assign grp_fu_397_p_din1 = grp_rayCast_fu_179_grp_fu_601_p_din1;

    assign grp_fu_397_p_opcode = grp_rayCast_fu_179_grp_fu_601_p_opcode;

    assign grp_fu_401_p_ce = grp_fu_597_ce;

    assign grp_fu_401_p_din0 = grp_fu_597_p0;

    assign grp_fu_401_p_din1 = grp_fu_597_p1;

    assign grp_fu_401_p_opcode = grp_fu_597_opcode;

    assign grp_fu_405_p_ce = grp_fu_605_ce;

    assign grp_fu_405_p_din0 = grp_fu_605_p0;

    assign grp_fu_405_p_din1 = grp_fu_605_p1;

    assign grp_fu_409_p_ce = grp_fu_609_ce;

    assign grp_fu_409_p_din0 = grp_fu_609_p0;

    assign grp_fu_409_p_din1 = grp_fu_609_p1;

    assign grp_fu_413_p_ce = grp_fu_620_ce;

    assign grp_fu_413_p_din0 = grp_fu_620_p0;

    assign grp_fu_413_p_din1 = grp_fu_620_p1;

    assign grp_fu_413_p_opcode = grp_fu_620_opcode;

    assign grp_fu_417_p_ce = grp_fu_646_ce;

    assign grp_fu_417_p_din0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din0;

    assign grp_fu_417_p_din1 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_grp_fu_646_p_din1;

    assign grp_rayCast_fu_179_ap_start = grp_rayCast_fu_179_ap_start_reg;

    assign grp_sin_or_cos_double_s_fu_421_p_din1 = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din1;

    assign grp_sin_or_cos_double_s_fu_421_p_din2 = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_624_p_din2;

    assign grp_sin_or_cos_double_s_fu_421_p_start = grp_sin_or_cos_double_s_fu_624_ap_start;

    assign grp_sin_or_cos_double_s_fu_432_p_din1 = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din1;

    assign grp_sin_or_cos_double_s_fu_432_p_din2 = grp_rayCast_fu_179_grp_sin_or_cos_double_s_fu_635_p_din2;

    assign grp_sin_or_cos_double_s_fu_432_p_start = grp_sin_or_cos_double_s_fu_635_ap_start;

    assign grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_ap_start_reg;

    assign icmp_ln162_fu_267_p2 = ((i_fu_96 == 9'd500) ? 1'b1 : 1'b0);

    assign icmp_ln168_fu_324_p2 = (($signed(d_reg_167) < $signed(33'd180)) ? 1'b1 : 1'b0);

    assign laserReading_address0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_address0;

    assign laserReading_ce0 = grp_updateSensor_Pipeline_VITIS_LOOP_173_3_fu_202_laserReading_ce0;

    assign mul_ln177_fu_253_p0 = mul_ln177_fu_253_p00;

    assign mul_ln177_fu_253_p00 = laserReading_offset;

    assign mul_ln177_fu_253_p1 = 18'd180;

    assign p_cast_fu_300_p4 = {{pf_q0[159:128]}};

    assign pf_d0 = {{bitcast_ln181_fu_418_p1}, {192'd0}};

    assign sext_ln168_fu_320_p1 = $signed(p_cast_fu_300_p4);

    assign theta_fu_296_p1 = grp_fu_239_p4;

    assign trunc_ln163_fu_284_p1 = pf_q1[63:0];

    assign trunc_ln205_fu_363_p1 = pf_q0[63:0];

    assign x_fu_288_p1 = trunc_ln163_fu_284_p1;

    assign y_fu_292_p1 = grp_fu_229_p4;

    assign zext_ln162_fu_279_p1 = i_fu_96;

    assign zext_ln168_fu_344_p1 = d_reg_167;

    always @(posedge ap_clk) begin
        pf_addr_3_reg_472[16:9] <= 8'b00000000;
    end

endmodule  //main_updateSensor
