/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_60_5_VITIS_LOOP_61_6_VITIS_LOOP_62_7 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    controlSequence_address0,
    controlSequence_ce0,
    controlSequence_we0,
    controlSequence_d0,
    controlSequence_address1,
    controlSequence_ce1,
    controlSequence_q1,
    mul3,
    grp_fu_242_p_din0,
    grp_fu_242_p_din1,
    grp_fu_242_p_opcode,
    grp_fu_242_p_dout0,
    grp_fu_242_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [4:0] controlSequence_address0;
    output controlSequence_ce0;
    output controlSequence_we0;
    output [31:0] controlSequence_d0;
    output [4:0] controlSequence_address1;
    output controlSequence_ce1;
    input [31:0] controlSequence_q1;
    input [31:0] mul3;
    output [31:0] grp_fu_242_p_din0;
    output [31:0] grp_fu_242_p_din1;
    output [0:0] grp_fu_242_p_opcode;
    input [31:0] grp_fu_242_p_dout0;
    output grp_fu_242_p_ce;

    reg ap_idle;
    reg controlSequence_ce0;
    reg controlSequence_we0;
    reg controlSequence_ce1;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln60_fu_118_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    wire   [1:0] select_ln61_fu_183_p3;
    reg   [1:0] select_ln61_reg_310;
    wire   [3:0] select_ln61_1_fu_191_p3;
    reg   [3:0] select_ln61_1_reg_315;
    wire   [2:0] empty_fu_199_p1;
    reg   [2:0] empty_reg_320;
    reg   [4:0] controlSequence_addr_reg_325;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter2_reg;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter3_reg;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter4_reg;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter5_reg;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter6_reg;
    reg   [4:0] controlSequence_addr_reg_325_pp0_iter7_reg;
    reg   [31:0] controlSequence_load_reg_331;
    reg   [31:0] sub4_reg_336;
    wire   [63:0] zext_ln63_fu_268_p1;
    wire    ap_block_pp0_stage0;
    reg   [1:0] dim_fu_52;
    wire   [1:0] add_ln62_fu_203_p2;
    wire    ap_loop_init;
    reg   [1:0] ap_sig_allocacmp_dim_load;
    reg   [3:0] i_fu_56;
    reg   [3:0] ap_sig_allocacmp_i_load;
    reg   [5:0] indvar_flatten_fu_60;
    wire   [5:0] select_ln61_2_fu_215_p3;
    reg   [5:0] ap_sig_allocacmp_indvar_flatten_load;
    reg   [11:0] indvar_flatten11_fu_64;
    wire   [11:0] add_ln60_fu_124_p2;
    reg   [11:0] ap_sig_allocacmp_indvar_flatten11_load;
    wire   [0:0] icmp_ln61_fu_139_p2;
    wire   [0:0] icmp_ln62_fu_159_p2;
    wire   [0:0] xor_ln60_fu_153_p2;
    wire   [3:0] select_ln60_fu_145_p3;
    wire   [0:0] and_ln60_fu_165_p2;
    wire   [0:0] or_ln61_fu_177_p2;
    wire   [3:0] add_ln61_fu_171_p2;
    wire   [5:0] add_ln61_1_fu_209_p2;
    wire   [4:0] p_shl3_fu_246_p3;
    wire   [4:0] zext_ln61_fu_243_p1;
    wire   [4:0] zext_ln62_fu_259_p1;
    wire   [4:0] empty_8_fu_253_p2;
    wire   [4:0] add_ln63_fu_262_p2;
    wire    ap_block_pp0_stage0_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 dim_fu_52 = 2'd0;
        #0 i_fu_56 = 4'd0;
        #0 indvar_flatten_fu_60 = 6'd0;
        #0 indvar_flatten11_fu_64 = 12'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter7_reg == 1'b1))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln60_fu_118_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                dim_fu_52 <= add_ln62_fu_203_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                dim_fu_52 <= 2'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln60_fu_118_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                i_fu_56 <= select_ln61_1_fu_191_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                i_fu_56 <= 4'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln60_fu_118_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                indvar_flatten11_fu_64 <= add_ln60_fu_124_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                indvar_flatten11_fu_64 <= 12'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln60_fu_118_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                indvar_flatten_fu_60 <= select_ln61_2_fu_215_p3;
            end else if ((ap_loop_init == 1'b1)) begin
                indvar_flatten_fu_60 <= 6'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
            controlSequence_addr_reg_325 <= zext_ln63_fu_268_p1;
            empty_reg_320 <= empty_fu_199_p1;
            select_ln61_1_reg_315 <= select_ln61_1_fu_191_p3;
            select_ln61_reg_310 <= select_ln61_fu_183_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
            controlSequence_addr_reg_325_pp0_iter2_reg <= controlSequence_addr_reg_325;
            controlSequence_addr_reg_325_pp0_iter3_reg <= controlSequence_addr_reg_325_pp0_iter2_reg;
            controlSequence_addr_reg_325_pp0_iter4_reg <= controlSequence_addr_reg_325_pp0_iter3_reg;
            controlSequence_addr_reg_325_pp0_iter5_reg <= controlSequence_addr_reg_325_pp0_iter4_reg;
            controlSequence_addr_reg_325_pp0_iter6_reg <= controlSequence_addr_reg_325_pp0_iter5_reg;
            controlSequence_addr_reg_325_pp0_iter7_reg <= controlSequence_addr_reg_325_pp0_iter6_reg;
            sub4_reg_336 <= grp_fu_242_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
            controlSequence_load_reg_331 <= controlSequence_q1;
        end
    end

    always @(*) begin
        if (((icmp_ln60_fu_118_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter7_reg == 1'b1))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            ap_sig_allocacmp_dim_load = 2'd0;
        end else begin
            ap_sig_allocacmp_dim_load = dim_fu_52;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            ap_sig_allocacmp_i_load = 4'd0;
        end else begin
            ap_sig_allocacmp_i_load = i_fu_56;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            ap_sig_allocacmp_indvar_flatten11_load = 12'd0;
        end else begin
            ap_sig_allocacmp_indvar_flatten11_load = indvar_flatten11_fu_64;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            ap_sig_allocacmp_indvar_flatten_load = 6'd0;
        end else begin
            ap_sig_allocacmp_indvar_flatten_load = indvar_flatten_fu_60;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter8 == 1'b1))) begin
            controlSequence_ce0 = 1'b1;
        end else begin
            controlSequence_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            controlSequence_ce1 = 1'b1;
        end else begin
            controlSequence_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter8 == 1'b1))) begin
            controlSequence_we0 = 1'b1;
        end else begin
            controlSequence_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln60_fu_124_p2 = (ap_sig_allocacmp_indvar_flatten11_load + 12'd1);

    assign add_ln61_1_fu_209_p2 = (ap_sig_allocacmp_indvar_flatten_load + 6'd1);

    assign add_ln61_fu_171_p2 = (select_ln60_fu_145_p3 + 4'd1);

    assign add_ln62_fu_203_p2 = (select_ln61_fu_183_p3 + 2'd1);

    assign add_ln63_fu_262_p2 = (zext_ln62_fu_259_p1 + empty_8_fu_253_p2);

    assign and_ln60_fu_165_p2 = (xor_ln60_fu_153_p2 & icmp_ln62_fu_159_p2);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign controlSequence_address0 = controlSequence_addr_reg_325_pp0_iter7_reg;

    assign controlSequence_address1 = zext_ln63_fu_268_p1;

    assign controlSequence_d0 = sub4_reg_336;

    assign empty_8_fu_253_p2 = (p_shl3_fu_246_p3 - zext_ln61_fu_243_p1);

    assign empty_fu_199_p1 = select_ln61_1_fu_191_p3[2:0];

    assign grp_fu_242_p_ce = 1'b1;

    assign grp_fu_242_p_din0 = controlSequence_load_reg_331;

    assign grp_fu_242_p_din1 = mul3;

    assign grp_fu_242_p_opcode = 2'd1;

    assign icmp_ln60_fu_118_p2 = ((ap_sig_allocacmp_indvar_flatten11_load == 12'd3000) ? 1'b1 : 1'b0);

    assign icmp_ln61_fu_139_p2 = ((ap_sig_allocacmp_indvar_flatten_load == 6'd30) ? 1'b1 : 1'b0);

    assign icmp_ln62_fu_159_p2 = ((ap_sig_allocacmp_dim_load == 2'd3) ? 1'b1 : 1'b0);

    assign or_ln61_fu_177_p2 = (icmp_ln61_fu_139_p2 | and_ln60_fu_165_p2);

    assign p_shl3_fu_246_p3 = {{empty_reg_320}, {2'd0}};

    assign select_ln60_fu_145_p3 = ((icmp_ln61_fu_139_p2[0:0] == 1'b1) ? 4'd0 : ap_sig_allocacmp_i_load);

    assign select_ln61_1_fu_191_p3 = ((and_ln60_fu_165_p2[0:0] == 1'b1) ? add_ln61_fu_171_p2 : select_ln60_fu_145_p3);

    assign select_ln61_2_fu_215_p3 = ((icmp_ln61_fu_139_p2[0:0] == 1'b1) ? 6'd1 : add_ln61_1_fu_209_p2);

    assign select_ln61_fu_183_p3 = ((or_ln61_fu_177_p2[0:0] == 1'b1) ? 2'd0 : ap_sig_allocacmp_dim_load);

    assign xor_ln60_fu_153_p2 = (icmp_ln61_fu_139_p2 ^ 1'd1);

    assign zext_ln61_fu_243_p1 = select_ln61_1_reg_315;

    assign zext_ln62_fu_259_p1 = select_ln61_reg_310;

    assign zext_ln63_fu_268_p1 = add_ln63_fu_262_p2;

endmodule  //main_main_Pipeline_VITIS_LOOP_60_5_VITIS_LOOP_61_6_VITIS_LOOP_62_7
