/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_sin_or_cos_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    t_in,
    do_cos,
    ap_return
);

    parameter ap_ST_fsm_state1 = 32'd1;
    parameter ap_ST_fsm_state2 = 32'd2;
    parameter ap_ST_fsm_state3 = 32'd4;
    parameter ap_ST_fsm_state4 = 32'd8;
    parameter ap_ST_fsm_state5 = 32'd16;
    parameter ap_ST_fsm_state6 = 32'd32;
    parameter ap_ST_fsm_state7 = 32'd64;
    parameter ap_ST_fsm_state8 = 32'd128;
    parameter ap_ST_fsm_state9 = 32'd256;
    parameter ap_ST_fsm_state10 = 32'd512;
    parameter ap_ST_fsm_state11 = 32'd1024;
    parameter ap_ST_fsm_state12 = 32'd2048;
    parameter ap_ST_fsm_state13 = 32'd4096;
    parameter ap_ST_fsm_state14 = 32'd8192;
    parameter ap_ST_fsm_state15 = 32'd16384;
    parameter ap_ST_fsm_state16 = 32'd32768;
    parameter ap_ST_fsm_state17 = 32'd65536;
    parameter ap_ST_fsm_state18 = 32'd131072;
    parameter ap_ST_fsm_state19 = 32'd262144;
    parameter ap_ST_fsm_state20 = 32'd524288;
    parameter ap_ST_fsm_state21 = 32'd1048576;
    parameter ap_ST_fsm_state22 = 32'd2097152;
    parameter ap_ST_fsm_state23 = 32'd4194304;
    parameter ap_ST_fsm_state24 = 32'd8388608;
    parameter ap_ST_fsm_state25 = 32'd16777216;
    parameter ap_ST_fsm_state26 = 32'd33554432;
    parameter ap_ST_fsm_state27 = 32'd67108864;
    parameter ap_ST_fsm_state28 = 32'd134217728;
    parameter ap_ST_fsm_state29 = 32'd268435456;
    parameter ap_ST_fsm_state30 = 32'd536870912;
    parameter ap_ST_fsm_state31 = 32'd1073741824;
    parameter ap_ST_fsm_state32 = 32'd2147483648;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] t_in;
    input [0:0] do_cos;
    output [63:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;

    (* fsm_encoding = "none" *) reg   [31:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire   [3:0] ref_4oPi_table_256_address0;
    reg    ref_4oPi_table_256_ce0;
    wire   [255:0] ref_4oPi_table_256_q0;
    wire   [7:0] fourth_order_double_sin_cos_K0_address0;
    reg    fourth_order_double_sin_cos_K0_ce0;
    wire   [58:0] fourth_order_double_sin_cos_K0_q0;
    wire   [7:0] fourth_order_double_sin_cos_K1_address0;
    reg    fourth_order_double_sin_cos_K1_ce0;
    wire   [51:0] fourth_order_double_sin_cos_K1_q0;
    wire   [7:0] fourth_order_double_sin_cos_K2_address0;
    reg    fourth_order_double_sin_cos_K2_ce0;
    wire   [43:0] fourth_order_double_sin_cos_K2_q0;
    wire   [7:0] fourth_order_double_sin_cos_K3_address0;
    reg    fourth_order_double_sin_cos_K3_ce0;
    wire   [32:0] fourth_order_double_sin_cos_K3_q0;
    wire   [7:0] fourth_order_double_sin_cos_K4_address0;
    reg    fourth_order_double_sin_cos_K4_ce0;
    wire   [24:0] fourth_order_double_sin_cos_K4_q0;
    reg   [0:0] din_sign_reg_1234;
    wire   [10:0] din_exp_fu_364_p4;
    reg   [10:0] din_exp_reg_1240;
    wire   [51:0] din_sig_fu_374_p1;
    reg   [51:0] din_sig_reg_1247;
    wire   [0:0] closepath_fu_378_p2;
    reg   [0:0] closepath_reg_1253;
    wire   [6:0] trunc_ln398_fu_413_p1;
    reg   [6:0] trunc_ln398_reg_1265;
    reg   [255:0] table_256_reg_1270;
    wire    ap_CS_fsm_state2;
    reg  signed [169:0] Med_reg_1275;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    wire   [0:0] icmp_ln271_1_fu_447_p2;
    reg   [0:0] icmp_ln271_1_reg_1285;
    wire   [169:0] grp_fu_348_p2;
    reg   [169:0] h_reg_1291;
    wire    ap_CS_fsm_state8;
    reg   [123:0] Mx_bits_reg_1296;
    reg   [2:0] k_reg_1302;
    wire   [2:0] k_1_fu_479_p3;
    reg   [2:0] k_1_reg_1307;
    wire    ap_CS_fsm_state9;
    wire   [123:0] Mx_bits_3_fu_501_p3;
    reg   [123:0] Mx_bits_3_reg_1313;
    wire   [6:0] Mx_zeros_fu_556_p1;
    reg   [6:0] Mx_zeros_reg_1318;
    reg   [62:0] Mx_reg_1324;
    wire    ap_CS_fsm_state10;
    wire   [10:0] Ex_1_fu_593_p2;
    reg   [10:0] Ex_1_reg_1331;
    reg   [0:0] tmp_16_reg_1337;
    wire   [10:0] sub_ln506_fu_607_p2;
    reg   [10:0] sub_ln506_reg_1343;
    wire   [0:0] icmp_ln271_fu_613_p2;
    reg   [0:0] icmp_ln271_reg_1348;
    wire   [0:0] icmp_ln282_fu_618_p2;
    reg   [0:0] icmp_ln282_reg_1354;
    reg   [6:0] tmp_17_reg_1361;
    wire    ap_CS_fsm_state11;
    wire   [55:0] B_fu_659_p1;
    reg   [55:0] B_reg_1366;
    reg   [48:0] B_trunc_reg_1371;
    wire   [97:0] zext_ln25_fu_673_p1;
    reg   [97:0] zext_ln25_reg_1376;
    wire    ap_CS_fsm_state12;
    wire    ap_CS_fsm_state15;
    wire   [0:0] cos_basis_fu_723_p3;
    reg   [0:0] cos_basis_reg_1388;
    wire   [63:0] zext_ln32_fu_746_p1;
    reg   [63:0] zext_ln32_reg_1395;
    reg   [48:0] B_squared_reg_1412;
    wire    ap_CS_fsm_state16;
    reg  signed [51:0] fourth_order_double_sin_cos_K1_load_reg_1418;
    reg  signed [43:0] fourth_order_double_sin_cos_K2_load_reg_1423;
    wire   [97:0] zext_ln25_1_fu_762_p1;
    wire    ap_CS_fsm_state17;
    wire    ap_CS_fsm_state20;
    reg   [58:0] t1_reg_1470;
    wire    ap_CS_fsm_state21;
    reg   [55:0] trunc_ln_reg_1475;
    reg   [47:0] trunc_ln2_reg_1480;
    reg   [41:0] tmp_11_reg_1485;
    reg   [32:0] fourth_order_double_sin_cos_K3_load_reg_1490;
    reg   [34:0] tmp_12_reg_1495;
    reg   [24:0] fourth_order_double_sin_cos_K4_load_reg_1500;
    wire    ap_CS_fsm_state22;
    wire   [63:0] add_ln37_1_fu_863_p2;
    reg   [63:0] add_ln37_1_reg_1525;
    reg   [28:0] lshr_ln_reg_1530;
    wire    ap_CS_fsm_state23;
    reg   [36:0] tmp_13_reg_1535;
    wire   [62:0] Mx_1_fu_889_p3;
    reg   [62:0] Mx_1_reg_1540;
    wire    ap_CS_fsm_state24;
    wire   [63:0] add_ln37_3_fu_906_p2;
    reg  signed [63:0] add_ln37_3_reg_1545;
    wire    ap_CS_fsm_state25;
    reg   [62:0] result_reg_1560;
    wire    ap_CS_fsm_state29;
    wire   [11:0] sub_ln252_fu_940_p2;
    reg   [11:0] sub_ln252_reg_1565;
    wire   [63:0] grp_scaled_fixed2ieee_63_1_s_fu_314_ap_return;
    reg   [63:0] resultf_reg_1570;
    wire    ap_CS_fsm_state31;
    wire    grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start;
    wire    grp_scaled_fixed2ieee_63_1_s_fu_314_ap_done;
    wire    grp_scaled_fixed2ieee_63_1_s_fu_314_ap_idle;
    wire    grp_scaled_fixed2ieee_63_1_s_fu_314_ap_ready;
    reg    grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg;
    wire    ap_CS_fsm_state30;
    wire   [63:0] zext_ln397_fu_408_p1;
    wire   [34:0] grp_fu_320_p0;
    wire   [24:0] grp_fu_320_p1;
    wire   [41:0] grp_fu_324_p0;
    wire   [32:0] grp_fu_324_p1;
    wire   [48:0] grp_fu_328_p0;
    reg   [48:0] grp_fu_332_p0;
    reg   [48:0] grp_fu_332_p1;
    wire   [48:0] grp_fu_336_p0;
    wire   [48:0] grp_fu_336_p1;
    wire   [55:0] grp_fu_340_p0;
    wire   [62:0] grp_fu_344_p1;
    wire   [52:0] grp_fu_348_p1;
    wire   [63:0] data_fu_352_p1;
    wire   [10:0] add_ln396_fu_384_p2;
    wire   [10:0] addr_fu_390_p3;
    wire   [3:0] tmp_s_fu_398_p4;
    wire   [255:0] zext_ln398_fu_417_p1;
    wire   [255:0] shl_ln398_fu_420_p2;
    wire   [52:0] X_fu_435_p3;
    wire   [0:0] tmp_fu_472_p3;
    wire   [0:0] xor_ln451_fu_485_p2;
    wire   [0:0] and_ln451_fu_490_p2;
    wire   [123:0] Mx_bits_1_fu_496_p2;
    wire   [60:0] tmp_24_fu_508_p4;
    wire   [61:0] t_fu_518_p3;
    reg   [61:0] tmp_6_fu_526_p4;
    wire   [62:0] tmp_7_fu_536_p3;
    wire  signed [63:0] sext_ln75_fu_544_p1;
    reg   [63:0] tmp_8_fu_548_p3;
    wire   [10:0] Ex_fu_560_p2;
    wire   [123:0] zext_ln504_fu_575_p1;
    wire   [123:0] shl_ln504_fu_578_p2;
    wire   [10:0] select_ln453_fu_565_p3;
    wire   [10:0] zext_ln505_fu_572_p1;
    wire   [10:0] select_ln506_fu_623_p3;
    wire   [62:0] zext_ln506_fu_628_p1;
    wire   [62:0] lshr_ln506_fu_632_p2;
    wire   [62:0] shl_ln506_fu_637_p2;
    wire   [62:0] x_1_fu_642_p3;
    wire   [0:0] tmp_9_fu_678_p17;
    wire   [0:0] tmp_9_fu_678_p19;
    wire   [0:0] xor_ln242_fu_717_p2;
    wire   [0:0] sin_basis_fu_731_p3;
    wire   [7:0] A_fu_739_p3;
    wire   [97:0] grp_fu_332_p2;
    wire   [107:0] grp_fu_340_p2;
    wire   [92:0] grp_fu_328_p2;
    wire   [97:0] grp_fu_336_p2;
    wire   [62:0] t1_1_fu_824_p3;
    wire  signed [63:0] sext_ln37_fu_847_p1;
    wire  signed [63:0] sext_ln37_1_fu_851_p1;
    wire   [63:0] add_ln37_fu_854_p2;
    wire  signed [63:0] sext_ln37_2_fu_860_p1;
    wire   [59:0] grp_fu_320_p2;
    wire   [74:0] grp_fu_324_p2;
    wire   [63:0] zext_ln37_2_fu_895_p1;
    wire   [63:0] add_ln37_2_fu_898_p2;
    wire   [63:0] zext_ln37_fu_903_p1;
    wire   [125:0] grp_fu_344_p2;
    wire   [10:0] Ex_2_fu_920_p3;
    wire  signed [11:0] sext_ln252_fu_936_p1;
    wire    ap_CS_fsm_state32;
    wire   [63:0] data_3_fu_946_p1;
    wire   [0:0] tmp_4_fu_977_p33;
    wire   [3:0] index_fu_971_p3;
    wire   [0:0] tmp_10_fu_1049_p33;
    wire   [0:0] tmp_4_fu_977_p35;
    wire   [0:0] tmp_10_fu_1049_p35;
    wire   [0:0] select_ln242_fu_1121_p3;
    wire   [0:0] results_sign_fu_949_p3;
    wire   [0:0] xor_ln278_fu_1138_p2;
    wire   [0:0] results_sign_1_fu_1128_p2;
    wire   [0:0] xor_ln282_fu_1155_p2;
    wire   [10:0] results_exp_fu_957_p4;
    wire   [0:0] and_ln271_fu_1134_p2;
    wire   [0:0] results_sign_3_fu_1143_p2;
    wire   [0:0] results_sign_4_fu_1160_p2;
    wire   [10:0] select_ln259_fu_1148_p3;
    wire   [10:0] results_exp_1_fu_1166_p3;
    wire   [0:0] and_ln271_1_fu_1189_p2;
    wire   [0:0] xor_ln271_fu_1193_p2;
    wire   [0:0] or_ln271_fu_1207_p2;
    wire   [51:0] select_ln271_fu_1199_p3;
    wire   [51:0] results_sig_fu_967_p1;
    wire   [0:0] results_sign_5_fu_1173_p3;
    wire   [10:0] results_exp_2_fu_1181_p3;
    wire   [51:0] results_sig_1_fu_1212_p3;
    wire   [63:0] t_4_fu_1220_p4;
    reg   [31:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    reg    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire   [59:0] grp_fu_320_p00;
    wire   [59:0] grp_fu_320_p10;
    wire   [74:0] grp_fu_324_p00;
    wire   [74:0] grp_fu_324_p10;
    wire   [92:0] grp_fu_328_p00;
    wire   [107:0] grp_fu_340_p00;
    wire   [125:0] grp_fu_344_p10;
    wire   [169:0] grp_fu_348_p10;
    wire   [2:0] tmp_9_fu_678_p1;
    wire   [2:0] tmp_9_fu_678_p3;
    wire   [2:0] tmp_9_fu_678_p5;
    wire   [2:0] tmp_9_fu_678_p7;
    wire  signed [2:0] tmp_9_fu_678_p9;
    wire  signed [2:0] tmp_9_fu_678_p11;
    wire  signed [2:0] tmp_9_fu_678_p13;
    wire  signed [2:0] tmp_9_fu_678_p15;
    wire   [3:0] tmp_4_fu_977_p1;
    wire   [3:0] tmp_4_fu_977_p3;
    wire   [3:0] tmp_4_fu_977_p5;
    wire   [3:0] tmp_4_fu_977_p7;
    wire   [3:0] tmp_4_fu_977_p9;
    wire   [3:0] tmp_4_fu_977_p11;
    wire   [3:0] tmp_4_fu_977_p13;
    wire   [3:0] tmp_4_fu_977_p15;
    wire  signed [3:0] tmp_4_fu_977_p17;
    wire  signed [3:0] tmp_4_fu_977_p19;
    wire  signed [3:0] tmp_4_fu_977_p21;
    wire  signed [3:0] tmp_4_fu_977_p23;
    wire  signed [3:0] tmp_4_fu_977_p25;
    wire  signed [3:0] tmp_4_fu_977_p27;
    wire  signed [3:0] tmp_4_fu_977_p29;
    wire  signed [3:0] tmp_4_fu_977_p31;
    wire   [3:0] tmp_10_fu_1049_p1;
    wire   [3:0] tmp_10_fu_1049_p3;
    wire   [3:0] tmp_10_fu_1049_p5;
    wire   [3:0] tmp_10_fu_1049_p7;
    wire   [3:0] tmp_10_fu_1049_p9;
    wire   [3:0] tmp_10_fu_1049_p11;
    wire   [3:0] tmp_10_fu_1049_p13;
    wire   [3:0] tmp_10_fu_1049_p15;
    wire  signed [3:0] tmp_10_fu_1049_p17;
    wire  signed [3:0] tmp_10_fu_1049_p19;
    wire  signed [3:0] tmp_10_fu_1049_p21;
    wire  signed [3:0] tmp_10_fu_1049_p23;
    wire  signed [3:0] tmp_10_fu_1049_p25;
    wire  signed [3:0] tmp_10_fu_1049_p27;
    wire  signed [3:0] tmp_10_fu_1049_p29;
    wire  signed [3:0] tmp_10_fu_1049_p31;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 32'd1;
        #0 grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg = 1'b0;
    end

    main_sin_or_cos_double_s_ref_4oPi_table_256_ROM_AUTO_1R #(
        .DataWidth(256),
        .AddressRange(10),
        .AddressWidth(4)
    ) ref_4oPi_table_256_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(ref_4oPi_table_256_address0),
        .ce0(ref_4oPi_table_256_ce0),
        .q0(ref_4oPi_table_256_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K0_ROM_1P_LUTRAM_1R #(
        .DataWidth(59),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K0_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K0_address0),
        .ce0(fourth_order_double_sin_cos_K0_ce0),
        .q0(fourth_order_double_sin_cos_K0_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K1_ROM_1P_LUTRAM_1R #(
        .DataWidth(52),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K1_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K1_address0),
        .ce0(fourth_order_double_sin_cos_K1_ce0),
        .q0(fourth_order_double_sin_cos_K1_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K2_ROM_1P_LUTRAM_1R #(
        .DataWidth(44),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K2_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K2_address0),
        .ce0(fourth_order_double_sin_cos_K2_ce0),
        .q0(fourth_order_double_sin_cos_K2_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K3_ROM_1P_LUTRAM_1R #(
        .DataWidth(33),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K3_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K3_address0),
        .ce0(fourth_order_double_sin_cos_K3_ce0),
        .q0(fourth_order_double_sin_cos_K3_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K4_ROM_1P_LUTRAM_1R #(
        .DataWidth(25),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K4_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K4_address0),
        .ce0(fourth_order_double_sin_cos_K4_ce0),
        .q0(fourth_order_double_sin_cos_K4_q0)
    );

    main_scaled_fixed2ieee_63_1_s grp_scaled_fixed2ieee_63_1_s_fu_314 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start),
        .ap_done(grp_scaled_fixed2ieee_63_1_s_fu_314_ap_done),
        .ap_idle(grp_scaled_fixed2ieee_63_1_s_fu_314_ap_idle),
        .ap_ready(grp_scaled_fixed2ieee_63_1_s_fu_314_ap_ready),
        .in_val(result_reg_1560),
        .prescale(sub_ln252_reg_1565),
        .ap_return(grp_scaled_fixed2ieee_63_1_s_fu_314_ap_return)
    );

    main_mul_35ns_25ns_60_2_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(35),
        .din1_WIDTH(25),
        .dout_WIDTH(60)
    ) mul_35ns_25ns_60_2_1_U55 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_320_p0),
        .din1(grp_fu_320_p1),
        .ce(1'b1),
        .dout(grp_fu_320_p2)
    );

    main_mul_42ns_33ns_75_2_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(42),
        .din1_WIDTH(33),
        .dout_WIDTH(75)
    ) mul_42ns_33ns_75_2_1_U56 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_324_p0),
        .din1(grp_fu_324_p1),
        .ce(1'b1),
        .dout(grp_fu_324_p2)
    );

    main_mul_49ns_44s_93_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(44),
        .dout_WIDTH(93)
    ) mul_49ns_44s_93_5_1_U57 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_328_p0),
        .din1(fourth_order_double_sin_cos_K2_load_reg_1423),
        .ce(1'b1),
        .dout(grp_fu_328_p2)
    );

    main_mul_49ns_49ns_98_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(49),
        .dout_WIDTH(98)
    ) mul_49ns_49ns_98_5_1_U58 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_332_p0),
        .din1(grp_fu_332_p1),
        .ce(1'b1),
        .dout(grp_fu_332_p2)
    );

    main_mul_49ns_49ns_98_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(49),
        .dout_WIDTH(98)
    ) mul_49ns_49ns_98_5_1_U59 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_336_p0),
        .din1(grp_fu_336_p1),
        .ce(1'b1),
        .dout(grp_fu_336_p2)
    );

    main_mul_56ns_52s_108_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(56),
        .din1_WIDTH(52),
        .dout_WIDTH(108)
    ) mul_56ns_52s_108_5_1_U60 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_340_p0),
        .din1(fourth_order_double_sin_cos_K1_load_reg_1418),
        .ce(1'b1),
        .dout(grp_fu_340_p2)
    );

    main_mul_64s_63ns_126_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(64),
        .din1_WIDTH(63),
        .dout_WIDTH(126)
    ) mul_64s_63ns_126_5_1_U61 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_ln37_3_reg_1545),
        .din1(grp_fu_344_p1),
        .ce(1'b1),
        .dout(grp_fu_344_p2)
    );

    main_mul_170s_53ns_170_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(170),
        .din1_WIDTH(53),
        .dout_WIDTH(170)
    ) mul_170s_53ns_170_5_1_U62 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(Med_reg_1275),
        .din1(grp_fu_348_p1),
        .ce(1'b1),
        .dout(grp_fu_348_p2)
    );

    main_sparsemux_17_3_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(3'h0),
        .din0_WIDTH(1),
        .CASE1(3'h1),
        .din1_WIDTH(1),
        .CASE2(3'h2),
        .din2_WIDTH(1),
        .CASE3(3'h3),
        .din3_WIDTH(1),
        .CASE4(3'h4),
        .din4_WIDTH(1),
        .CASE5(3'h5),
        .din5_WIDTH(1),
        .CASE6(3'h6),
        .din6_WIDTH(1),
        .CASE7(3'h7),
        .din7_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(3),
        .dout_WIDTH(1)
    ) sparsemux_17_3_1_1_1_U63 (
        .din0(1'd0),
        .din1(1'd1),
        .din2(1'd1),
        .din3(1'd0),
        .din4(1'd0),
        .din5(1'd1),
        .din6(1'd1),
        .din7(1'd0),
        .def (tmp_9_fu_678_p17),
        .sel (k_1_reg_1307),
        .dout(tmp_9_fu_678_p19)
    );

    main_sparsemux_33_4_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(4'h0),
        .din0_WIDTH(1),
        .CASE1(4'h1),
        .din1_WIDTH(1),
        .CASE2(4'h2),
        .din2_WIDTH(1),
        .CASE3(4'h3),
        .din3_WIDTH(1),
        .CASE4(4'h4),
        .din4_WIDTH(1),
        .CASE5(4'h5),
        .din5_WIDTH(1),
        .CASE6(4'h6),
        .din6_WIDTH(1),
        .CASE7(4'h7),
        .din7_WIDTH(1),
        .CASE8(4'h8),
        .din8_WIDTH(1),
        .CASE9(4'h9),
        .din9_WIDTH(1),
        .CASE10(4'hA),
        .din10_WIDTH(1),
        .CASE11(4'hB),
        .din11_WIDTH(1),
        .CASE12(4'hC),
        .din12_WIDTH(1),
        .CASE13(4'hD),
        .din13_WIDTH(1),
        .CASE14(4'hE),
        .din14_WIDTH(1),
        .CASE15(4'hF),
        .din15_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(4),
        .dout_WIDTH(1)
    ) sparsemux_33_4_1_1_1_U64 (
        .din0 (1'd0),
        .din1 (1'd0),
        .din2 (1'd0),
        .din3 (1'd1),
        .din4 (1'd1),
        .din5 (1'd1),
        .din6 (1'd1),
        .din7 (1'd0),
        .din8 (1'd0),
        .din9 (1'd1),
        .din10(1'd1),
        .din11(1'd1),
        .din12(1'd1),
        .din13(1'd0),
        .din14(1'd0),
        .din15(1'd0),
        .def  (tmp_4_fu_977_p33),
        .sel  (index_fu_971_p3),
        .dout (tmp_4_fu_977_p35)
    );

    main_sparsemux_33_4_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(4'h0),
        .din0_WIDTH(1),
        .CASE1(4'h1),
        .din1_WIDTH(1),
        .CASE2(4'h2),
        .din2_WIDTH(1),
        .CASE3(4'h3),
        .din3_WIDTH(1),
        .CASE4(4'h4),
        .din4_WIDTH(1),
        .CASE5(4'h5),
        .din5_WIDTH(1),
        .CASE6(4'h6),
        .din6_WIDTH(1),
        .CASE7(4'h7),
        .din7_WIDTH(1),
        .CASE8(4'h8),
        .din8_WIDTH(1),
        .CASE9(4'h9),
        .din9_WIDTH(1),
        .CASE10(4'hA),
        .din10_WIDTH(1),
        .CASE11(4'hB),
        .din11_WIDTH(1),
        .CASE12(4'hC),
        .din12_WIDTH(1),
        .CASE13(4'hD),
        .din13_WIDTH(1),
        .CASE14(4'hE),
        .din14_WIDTH(1),
        .CASE15(4'hF),
        .din15_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(4),
        .dout_WIDTH(1)
    ) sparsemux_33_4_1_1_1_U65 (
        .din0 (1'd0),
        .din1 (1'd0),
        .din2 (1'd1),
        .din3 (1'd0),
        .din4 (1'd1),
        .din5 (1'd1),
        .din6 (1'd0),
        .din7 (1'd1),
        .din8 (1'd1),
        .din9 (1'd0),
        .din10(1'd1),
        .din11(1'd1),
        .din12(1'd0),
        .din13(1'd1),
        .din14(1'd0),
        .din15(1'd0),
        .def  (tmp_10_fu_1049_p33),
        .sel  (index_fu_971_p3),
        .dout (tmp_10_fu_1049_p35)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state30)) begin
                grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg <= 1'b1;
            end else if ((grp_scaled_fixed2ieee_63_1_s_fu_314_ap_ready == 1'b1)) begin
                grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            B_reg_1366 <= B_fu_659_p1;
            B_trunc_reg_1371 <= {{x_1_fu_642_p3[55:7]}};
            tmp_17_reg_1361 <= {{x_1_fu_642_p3[62:56]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state16)) begin
            B_squared_reg_1412 <= {{grp_fu_332_p2[97:49]}};
            fourth_order_double_sin_cos_K1_load_reg_1418 <= fourth_order_double_sin_cos_K1_q0;
            fourth_order_double_sin_cos_K2_load_reg_1423 <= fourth_order_double_sin_cos_K2_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            Ex_1_reg_1331 <= Ex_1_fu_593_p2;
            Mx_reg_1324 <= {{shl_ln504_fu_578_p2[123:61]}};
            icmp_ln271_reg_1348 <= icmp_ln271_fu_613_p2;
            icmp_ln282_reg_1354 <= icmp_ln282_fu_618_p2;
            sub_ln506_reg_1343 <= sub_ln506_fu_607_p2;
            tmp_16_reg_1337 <= Ex_1_fu_593_p2[32'd10];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            Med_reg_1275 <= {{shl_ln398_fu_420_p2[255:86]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state24)) begin
            Mx_1_reg_1540 <= Mx_1_fu_889_p3;
            add_ln37_3_reg_1545 <= add_ln37_3_fu_906_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            Mx_bits_3_reg_1313 <= Mx_bits_3_fu_501_p3;
            Mx_zeros_reg_1318 <= Mx_zeros_fu_556_p1;
            k_1_reg_1307 <= k_1_fu_479_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            Mx_bits_reg_1296 <= {{grp_fu_348_p2[166:43]}};
            h_reg_1291 <= grp_fu_348_p2;
            k_reg_1302 <= {{grp_fu_348_p2[169:167]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state22)) begin
            add_ln37_1_reg_1525 <= add_ln37_1_fu_863_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            closepath_reg_1253 <= closepath_fu_378_p2;
            din_exp_reg_1240 <= {{data_fu_352_p1[62:52]}};
            din_sig_reg_1247 <= din_sig_fu_374_p1;
            din_sign_reg_1234 <= data_fu_352_p1[32'd63];
            trunc_ln398_reg_1265 <= trunc_ln398_fu_413_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            cos_basis_reg_1388 <= cos_basis_fu_723_p3;
            zext_ln32_reg_1395[7 : 0] <= zext_ln32_fu_746_p1[7 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state21)) begin
            fourth_order_double_sin_cos_K3_load_reg_1490 <= fourth_order_double_sin_cos_K3_q0;
            fourth_order_double_sin_cos_K4_load_reg_1500 <= fourth_order_double_sin_cos_K4_q0;
            t1_reg_1470 <= fourth_order_double_sin_cos_K0_q0;
            tmp_11_reg_1485 <= {{grp_fu_332_p2[97:56]}};
            tmp_12_reg_1495 <= {{grp_fu_336_p2[97:63]}};
            trunc_ln2_reg_1480 <= {{grp_fu_328_p2[92:45]}};
            trunc_ln_reg_1475 <= {{grp_fu_340_p2[107:52]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            icmp_ln271_1_reg_1285 <= icmp_ln271_1_fu_447_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state23)) begin
            lshr_ln_reg_1530 <= {{grp_fu_320_p2[59:31]}};
            tmp_13_reg_1535  <= {{grp_fu_324_p2[74:38]}};
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state29)) begin
            result_reg_1560 <= {{grp_fu_344_p2[125:63]}};
            sub_ln252_reg_1565 <= sub_ln252_fu_940_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state31)) begin
            resultf_reg_1570 <= grp_scaled_fixed2ieee_63_1_s_fu_314_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            table_256_reg_1270 <= ref_4oPi_table_256_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            zext_ln25_reg_1376[48 : 0] <= zext_ln25_fu_673_p1[48 : 0];
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    always @(*) begin
        if ((grp_scaled_fixed2ieee_63_1_s_fu_314_ap_done == 1'b0)) begin
            ap_ST_fsm_state31_blk = 1'b1;
        end else begin
            ap_ST_fsm_state31_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state32) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state32)) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state20)) begin
            fourth_order_double_sin_cos_K0_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            fourth_order_double_sin_cos_K1_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            fourth_order_double_sin_cos_K2_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state20)) begin
            fourth_order_double_sin_cos_K3_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state20)) begin
            fourth_order_double_sin_cos_K4_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K4_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_332_p0 = zext_ln25_1_fu_762_p1;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_332_p0 = zext_ln25_fu_673_p1;
        end else begin
            grp_fu_332_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            grp_fu_332_p1 = zext_ln25_reg_1376;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_332_p1 = zext_ln25_fu_673_p1;
        end else begin
            grp_fu_332_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ref_4oPi_table_256_ce0 = 1'b1;
        end else begin
            ref_4oPi_table_256_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                if (((grp_scaled_fixed2ieee_63_1_s_fu_314_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state31))) begin
                    ap_NS_fsm = ap_ST_fsm_state32;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state31;
                end
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign A_fu_739_p3 = {{sin_basis_fu_731_p3}, {tmp_17_reg_1361}};

    assign B_fu_659_p1 = x_1_fu_642_p3[55:0];

    assign Ex_1_fu_593_p2 = (select_ln453_fu_565_p3 - zext_ln505_fu_572_p1);

    assign Ex_2_fu_920_p3 = ((cos_basis_reg_1388[0:0] == 1'b1) ? 11'd0 : Ex_1_reg_1331);

    assign Ex_fu_560_p2 = ($signed(din_exp_reg_1240) + $signed(11'd1027));

    assign Mx_1_fu_889_p3 = ((cos_basis_reg_1388[0:0] == 1'b1) ? 63'd9223372036854775807 : Mx_reg_1324);

    assign Mx_bits_1_fu_496_p2 = (124'd0 - Mx_bits_reg_1296);

    assign Mx_bits_3_fu_501_p3 = ((and_ln451_fu_490_p2[0:0] == 1'b1) ? Mx_bits_1_fu_496_p2 : Mx_bits_reg_1296);

    assign Mx_zeros_fu_556_p1 = tmp_8_fu_548_p3[6:0];

    assign X_fu_435_p3 = {{1'd1}, {din_sig_reg_1247}};

    assign add_ln37_1_fu_863_p2 = ($signed(add_ln37_fu_854_p2) + $signed(sext_ln37_2_fu_860_p1));

    assign add_ln37_2_fu_898_p2 = (add_ln37_1_reg_1525 + zext_ln37_2_fu_895_p1);

    assign add_ln37_3_fu_906_p2 = (add_ln37_2_fu_898_p2 + zext_ln37_fu_903_p1);

    assign add_ln37_fu_854_p2 = ($signed(sext_ln37_fu_847_p1) + $signed(sext_ln37_1_fu_851_p1));

    assign add_ln396_fu_384_p2 = ($signed(din_exp_fu_364_p4) + $signed(11'd1101));

    assign addr_fu_390_p3 = ((closepath_fu_378_p2[0:0] == 1'b1) ? 11'd74 : add_ln396_fu_384_p2);

    assign and_ln271_1_fu_1189_p2 = (icmp_ln271_reg_1348 & icmp_ln271_1_reg_1285);

    assign and_ln271_fu_1134_p2 = (icmp_ln271_reg_1348 & icmp_ln271_1_reg_1285);

    assign and_ln451_fu_490_p2 = (xor_ln451_fu_485_p2 & tmp_fu_472_p3);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];

    assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];

    assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];

    assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];

    assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign ap_return = t_4_fu_1220_p4;

    assign closepath_fu_378_p2 = ((din_exp_fu_364_p4 < 11'd1022) ? 1'b1 : 1'b0);

    assign cos_basis_fu_723_p3 = ((do_cos[0:0] == 1'b1) ? xor_ln242_fu_717_p2 : tmp_9_fu_678_p19);

    assign data_3_fu_946_p1 = resultf_reg_1570;

    assign data_fu_352_p1 = t_in;

    assign din_exp_fu_364_p4 = {{data_fu_352_p1[62:52]}};

    assign din_sig_fu_374_p1 = data_fu_352_p1[51:0];

    assign fourth_order_double_sin_cos_K0_address0 = zext_ln32_reg_1395;

    assign fourth_order_double_sin_cos_K1_address0 = zext_ln32_fu_746_p1;

    assign fourth_order_double_sin_cos_K2_address0 = zext_ln32_fu_746_p1;

    assign fourth_order_double_sin_cos_K3_address0 = zext_ln32_reg_1395;

    assign fourth_order_double_sin_cos_K4_address0 = zext_ln32_reg_1395;

    assign grp_fu_320_p0 = grp_fu_320_p00;

    assign grp_fu_320_p00 = tmp_12_reg_1495;

    assign grp_fu_320_p1 = grp_fu_320_p10;

    assign grp_fu_320_p10 = fourth_order_double_sin_cos_K4_load_reg_1500;

    assign grp_fu_324_p0 = grp_fu_324_p00;

    assign grp_fu_324_p00 = tmp_11_reg_1485;

    assign grp_fu_324_p1 = grp_fu_324_p10;

    assign grp_fu_324_p10 = fourth_order_double_sin_cos_K3_load_reg_1490;

    assign grp_fu_328_p0 = grp_fu_328_p00;

    assign grp_fu_328_p00 = B_squared_reg_1412;

    assign grp_fu_336_p0 = zext_ln25_1_fu_762_p1;

    assign grp_fu_336_p1 = zext_ln25_1_fu_762_p1;

    assign grp_fu_340_p0 = grp_fu_340_p00;

    assign grp_fu_340_p00 = B_reg_1366;

    assign grp_fu_344_p1 = grp_fu_344_p10;

    assign grp_fu_344_p10 = Mx_1_reg_1540;

    assign grp_fu_348_p1 = grp_fu_348_p10;

    assign grp_fu_348_p10 = X_fu_435_p3;

    assign grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start = grp_scaled_fixed2ieee_63_1_s_fu_314_ap_start_reg;

    assign icmp_ln271_1_fu_447_p2 = ((din_sig_reg_1247 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln271_fu_613_p2 = ((din_exp_reg_1240 == 11'd0) ? 1'b1 : 1'b0);

    assign icmp_ln282_fu_618_p2 = ((din_exp_reg_1240 == 11'd2047) ? 1'b1 : 1'b0);

    assign index_fu_971_p3 = {{din_sign_reg_1234}, {k_1_reg_1307}};

    assign k_1_fu_479_p3 = ((closepath_reg_1253[0:0] == 1'b1) ? 3'd0 : k_reg_1302);

    assign lshr_ln506_fu_632_p2 = Mx_reg_1324 >> zext_ln506_fu_628_p1;

    assign or_ln271_fu_1207_p2 = (icmp_ln282_reg_1354 | and_ln271_fu_1134_p2);

    assign ref_4oPi_table_256_address0 = zext_ln397_fu_408_p1;

    assign results_exp_1_fu_1166_p3 = ((icmp_ln282_reg_1354[0:0] == 1'b1) ? 11'd2047 : results_exp_fu_957_p4);

    assign results_exp_2_fu_1181_p3 = ((and_ln271_fu_1134_p2[0:0] == 1'b1) ? select_ln259_fu_1148_p3 : results_exp_1_fu_1166_p3);

    assign results_exp_fu_957_p4 = {{data_3_fu_946_p1[62:52]}};

    assign results_sig_1_fu_1212_p3 = ((or_ln271_fu_1207_p2[0:0] == 1'b1) ? select_ln271_fu_1199_p3 : results_sig_fu_967_p1);

    assign results_sig_fu_967_p1 = data_3_fu_946_p1[51:0];

    assign results_sign_1_fu_1128_p2 = (select_ln242_fu_1121_p3 | results_sign_fu_949_p3);

    assign results_sign_3_fu_1143_p2 = (xor_ln278_fu_1138_p2 & din_sign_reg_1234);

    assign results_sign_4_fu_1160_p2 = (xor_ln282_fu_1155_p2 & results_sign_1_fu_1128_p2);

    assign results_sign_5_fu_1173_p3 = ((and_ln271_fu_1134_p2[0:0] == 1'b1) ? results_sign_3_fu_1143_p2 : results_sign_4_fu_1160_p2);

    assign results_sign_fu_949_p3 = data_3_fu_946_p1[32'd63];

    assign select_ln242_fu_1121_p3 = ((cos_basis_reg_1388[0:0] == 1'b1) ? tmp_4_fu_977_p35 : tmp_10_fu_1049_p35);

    assign select_ln259_fu_1148_p3 = ((do_cos[0:0] == 1'b1) ? 11'd1023 : 11'd0);

    assign select_ln271_fu_1199_p3 = ((xor_ln271_fu_1193_p2[0:0] == 1'b1) ? 52'd4503599627370495 : 52'd0);

    assign select_ln453_fu_565_p3 = ((closepath_reg_1253[0:0] == 1'b1) ? Ex_fu_560_p2 : 11'd0);

    assign select_ln506_fu_623_p3 = ((tmp_16_reg_1337[0:0] == 1'b1) ? sub_ln506_reg_1343 : Ex_1_reg_1331);

    assign sext_ln252_fu_936_p1 = $signed(Ex_2_fu_920_p3);

    assign sext_ln37_1_fu_851_p1 = $signed(trunc_ln_reg_1475);

    assign sext_ln37_2_fu_860_p1 = $signed(trunc_ln2_reg_1480);

    assign sext_ln37_fu_847_p1 = $signed(t1_1_fu_824_p3);

    assign sext_ln75_fu_544_p1 = $signed(tmp_7_fu_536_p3);

    assign shl_ln398_fu_420_p2 = table_256_reg_1270 << zext_ln398_fu_417_p1;

    assign shl_ln504_fu_578_p2 = Mx_bits_3_reg_1313 << zext_ln504_fu_575_p1;

    assign shl_ln506_fu_637_p2 = Mx_reg_1324 << zext_ln506_fu_628_p1;

    assign sin_basis_fu_731_p3 = ((do_cos[0:0] == 1'b1) ? tmp_9_fu_678_p19 : xor_ln242_fu_717_p2);

    assign sub_ln252_fu_940_p2 = ($signed(12'd0) - $signed(sext_ln252_fu_936_p1));

    assign sub_ln506_fu_607_p2 = (11'd0 - Ex_1_fu_593_p2);

    assign t1_1_fu_824_p3 = {{t1_reg_1470}, {4'd0}};

    assign t_4_fu_1220_p4 = {
        {{results_sign_5_fu_1173_p3}, {results_exp_2_fu_1181_p3}}, {results_sig_1_fu_1212_p3}
    };

    assign t_fu_518_p3 = {{tmp_24_fu_508_p4}, {1'd1}};

    assign tmp_10_fu_1049_p33 = 'bx;

    assign tmp_24_fu_508_p4 = {{Mx_bits_3_fu_501_p3[123:63]}};

    assign tmp_4_fu_977_p33 = 'bx;

    integer ap_tvar_int_0;

    always @(t_fu_518_p3) begin
        for (ap_tvar_int_0 = 62 - 1; ap_tvar_int_0 >= 0; ap_tvar_int_0 = ap_tvar_int_0 - 1) begin
            if (ap_tvar_int_0 > 61 - 0) begin
                tmp_6_fu_526_p4[ap_tvar_int_0] = 1'b0;
            end else begin
                tmp_6_fu_526_p4[ap_tvar_int_0] = t_fu_518_p3[61-ap_tvar_int_0];
            end
        end
    end

    assign tmp_7_fu_536_p3 = {{1'd1}, {tmp_6_fu_526_p4}};


    always @(sext_ln75_fu_544_p1) begin
        if (sext_ln75_fu_544_p1[0] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd0;
        end else if (sext_ln75_fu_544_p1[1] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd1;
        end else if (sext_ln75_fu_544_p1[2] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd2;
        end else if (sext_ln75_fu_544_p1[3] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd3;
        end else if (sext_ln75_fu_544_p1[4] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd4;
        end else if (sext_ln75_fu_544_p1[5] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd5;
        end else if (sext_ln75_fu_544_p1[6] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd6;
        end else if (sext_ln75_fu_544_p1[7] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd7;
        end else if (sext_ln75_fu_544_p1[8] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd8;
        end else if (sext_ln75_fu_544_p1[9] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd9;
        end else if (sext_ln75_fu_544_p1[10] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd10;
        end else if (sext_ln75_fu_544_p1[11] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd11;
        end else if (sext_ln75_fu_544_p1[12] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd12;
        end else if (sext_ln75_fu_544_p1[13] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd13;
        end else if (sext_ln75_fu_544_p1[14] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd14;
        end else if (sext_ln75_fu_544_p1[15] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd15;
        end else if (sext_ln75_fu_544_p1[16] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd16;
        end else if (sext_ln75_fu_544_p1[17] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd17;
        end else if (sext_ln75_fu_544_p1[18] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd18;
        end else if (sext_ln75_fu_544_p1[19] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd19;
        end else if (sext_ln75_fu_544_p1[20] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd20;
        end else if (sext_ln75_fu_544_p1[21] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd21;
        end else if (sext_ln75_fu_544_p1[22] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd22;
        end else if (sext_ln75_fu_544_p1[23] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd23;
        end else if (sext_ln75_fu_544_p1[24] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd24;
        end else if (sext_ln75_fu_544_p1[25] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd25;
        end else if (sext_ln75_fu_544_p1[26] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd26;
        end else if (sext_ln75_fu_544_p1[27] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd27;
        end else if (sext_ln75_fu_544_p1[28] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd28;
        end else if (sext_ln75_fu_544_p1[29] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd29;
        end else if (sext_ln75_fu_544_p1[30] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd30;
        end else if (sext_ln75_fu_544_p1[31] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd31;
        end else if (sext_ln75_fu_544_p1[32] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd32;
        end else if (sext_ln75_fu_544_p1[33] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd33;
        end else if (sext_ln75_fu_544_p1[34] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd34;
        end else if (sext_ln75_fu_544_p1[35] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd35;
        end else if (sext_ln75_fu_544_p1[36] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd36;
        end else if (sext_ln75_fu_544_p1[37] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd37;
        end else if (sext_ln75_fu_544_p1[38] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd38;
        end else if (sext_ln75_fu_544_p1[39] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd39;
        end else if (sext_ln75_fu_544_p1[40] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd40;
        end else if (sext_ln75_fu_544_p1[41] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd41;
        end else if (sext_ln75_fu_544_p1[42] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd42;
        end else if (sext_ln75_fu_544_p1[43] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd43;
        end else if (sext_ln75_fu_544_p1[44] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd44;
        end else if (sext_ln75_fu_544_p1[45] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd45;
        end else if (sext_ln75_fu_544_p1[46] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd46;
        end else if (sext_ln75_fu_544_p1[47] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd47;
        end else if (sext_ln75_fu_544_p1[48] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd48;
        end else if (sext_ln75_fu_544_p1[49] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd49;
        end else if (sext_ln75_fu_544_p1[50] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd50;
        end else if (sext_ln75_fu_544_p1[51] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd51;
        end else if (sext_ln75_fu_544_p1[52] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd52;
        end else if (sext_ln75_fu_544_p1[53] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd53;
        end else if (sext_ln75_fu_544_p1[54] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd54;
        end else if (sext_ln75_fu_544_p1[55] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd55;
        end else if (sext_ln75_fu_544_p1[56] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd56;
        end else if (sext_ln75_fu_544_p1[57] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd57;
        end else if (sext_ln75_fu_544_p1[58] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd58;
        end else if (sext_ln75_fu_544_p1[59] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd59;
        end else if (sext_ln75_fu_544_p1[60] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd60;
        end else if (sext_ln75_fu_544_p1[61] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd61;
        end else if (sext_ln75_fu_544_p1[62] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd62;
        end else if (sext_ln75_fu_544_p1[63] == 1'b1) begin
            tmp_8_fu_548_p3 = 64'd63;
        end else begin
            tmp_8_fu_548_p3 = 64'd64;
        end
    end

    assign tmp_9_fu_678_p17 = 'bx;

    assign tmp_fu_472_p3 = h_reg_1291[32'd167];

    assign tmp_s_fu_398_p4 = {{addr_fu_390_p3[10:7]}};

    assign trunc_ln398_fu_413_p1 = addr_fu_390_p3[6:0];

    assign x_1_fu_642_p3 = ((tmp_16_reg_1337[0:0] == 1'b1) ? lshr_ln506_fu_632_p2 : shl_ln506_fu_637_p2);

    assign xor_ln242_fu_717_p2 = (tmp_9_fu_678_p19 ^ 1'd1);

    assign xor_ln271_fu_1193_p2 = (1'd1 ^ and_ln271_1_fu_1189_p2);

    assign xor_ln278_fu_1138_p2 = (do_cos ^ 1'd1);

    assign xor_ln282_fu_1155_p2 = (icmp_ln282_reg_1354 ^ 1'd1);

    assign xor_ln451_fu_485_p2 = (closepath_reg_1253 ^ 1'd1);

    assign zext_ln25_1_fu_762_p1 = B_squared_reg_1412;

    assign zext_ln25_fu_673_p1 = B_trunc_reg_1371;

    assign zext_ln32_fu_746_p1 = A_fu_739_p3;

    assign zext_ln37_2_fu_895_p1 = tmp_13_reg_1535;

    assign zext_ln37_fu_903_p1 = lshr_ln_reg_1530;

    assign zext_ln397_fu_408_p1 = tmp_s_fu_398_p4;

    assign zext_ln398_fu_417_p1 = trunc_ln398_reg_1265;

    assign zext_ln504_fu_575_p1 = Mx_zeros_reg_1318;

    assign zext_ln505_fu_572_p1 = Mx_zeros_reg_1318;

    assign zext_ln506_fu_628_p1 = select_ln506_fu_623_p3;

    always @(posedge ap_clk) begin
        zext_ln25_reg_1376[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1395[63:8]  <= 56'b00000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_sin_or_cos_double_s
