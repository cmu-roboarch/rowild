/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_planRRT (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    this_0_0_0_0_address0,
    this_0_0_0_0_ce0,
    this_0_0_0_0_q0,
    this_0_0_0_1_address0,
    this_0_0_0_1_ce0,
    this_0_0_0_1_q0,
    this_0_0_0_2_address0,
    this_0_0_0_2_ce0,
    this_0_0_0_2_q0,
    this_0_0_1_0_address0,
    this_0_0_1_0_ce0,
    this_0_0_1_0_q0,
    this_0_0_1_1_address0,
    this_0_0_1_1_ce0,
    this_0_0_1_1_q0,
    this_0_0_1_2_address0,
    this_0_0_1_2_ce0,
    this_0_0_1_2_q0,
    this_0_0_2_0_address0,
    this_0_0_2_0_ce0,
    this_0_0_2_0_q0,
    this_0_0_2_1_address0,
    this_0_0_2_1_ce0,
    this_0_0_2_1_q0,
    this_0_0_2_2_address0,
    this_0_0_2_2_ce0,
    this_0_0_2_2_q0,
    this_0_0_3_0_address0,
    this_0_0_3_0_ce0,
    this_0_0_3_0_q0,
    this_0_0_3_1_address0,
    this_0_0_3_1_ce0,
    this_0_0_3_1_q0,
    this_0_0_3_2_address0,
    this_0_0_3_2_ce0,
    this_0_0_3_2_q0,
    this_0_0_4_0_address0,
    this_0_0_4_0_ce0,
    this_0_0_4_0_q0,
    this_0_0_4_1_address0,
    this_0_0_4_1_ce0,
    this_0_0_4_1_q0,
    this_0_0_4_2_address0,
    this_0_0_4_2_ce0,
    this_0_0_4_2_q0,
    this_0_0_5_0_address0,
    this_0_0_5_0_ce0,
    this_0_0_5_0_q0,
    this_0_0_5_1_address0,
    this_0_0_5_1_ce0,
    this_0_0_5_1_q0,
    this_0_0_5_2_address0,
    this_0_0_5_2_ce0,
    this_0_0_5_2_q0,
    this_0_0_6_0_address0,
    this_0_0_6_0_ce0,
    this_0_0_6_0_q0,
    this_0_0_6_1_address0,
    this_0_0_6_1_ce0,
    this_0_0_6_1_q0,
    this_0_0_6_2_address0,
    this_0_0_6_2_ce0,
    this_0_0_6_2_q0,
    this_0_0_7_0_address0,
    this_0_0_7_0_ce0,
    this_0_0_7_0_q0,
    this_0_0_7_1_address0,
    this_0_0_7_1_ce0,
    this_0_0_7_1_q0,
    this_0_0_7_2_address0,
    this_0_0_7_2_ce0,
    this_0_0_7_2_q0,
    this_0_0_8_0_address0,
    this_0_0_8_0_ce0,
    this_0_0_8_0_q0,
    this_0_0_8_1_address0,
    this_0_0_8_1_ce0,
    this_0_0_8_1_q0,
    this_0_0_8_2_address0,
    this_0_0_8_2_ce0,
    this_0_0_8_2_q0,
    this_0_1_address0,
    this_0_1_ce0,
    this_0_1_q0,
    this_0_1_address1,
    this_0_1_ce1,
    this_0_1_q1,
    this_4_0_0_address0,
    this_4_0_0_ce0,
    this_4_0_0_q0,
    this_4_0_1_address0,
    this_4_0_1_ce0,
    this_4_0_1_q0,
    this_4_0_2_address0,
    this_4_0_2_ce0,
    this_4_0_2_q0,
    this_4_0_3_address0,
    this_4_0_3_ce0,
    this_4_0_3_q0,
    this_4_1_0_address0,
    this_4_1_0_ce0,
    this_4_1_0_q0,
    this_4_1_1_address0,
    this_4_1_1_ce0,
    this_4_1_1_q0,
    this_4_1_2_address0,
    this_4_1_2_ce0,
    this_4_1_2_q0,
    this_4_1_3_address0,
    this_4_1_3_ce0,
    this_4_1_3_q0,
    this_4_2_0_address0,
    this_4_2_0_ce0,
    this_4_2_0_q0,
    this_4_2_1_address0,
    this_4_2_1_ce0,
    this_4_2_1_q0,
    this_4_2_2_address0,
    this_4_2_2_ce0,
    this_4_2_2_q0,
    this_4_2_3_address0,
    this_4_2_3_ce0,
    this_4_2_3_q0,
    this_4_3_0_address0,
    this_4_3_0_ce0,
    this_4_3_0_q0,
    this_4_3_1_address0,
    this_4_3_1_ce0,
    this_4_3_1_q0,
    this_4_3_2_address0,
    this_4_3_2_ce0,
    this_4_3_2_q0,
    this_4_3_3_address0,
    this_4_3_3_ce0,
    this_4_3_3_q0,
    this_5_0_0_address0,
    this_5_0_0_ce0,
    this_5_0_0_we0,
    this_5_0_0_d0,
    this_5_0_0_q0,
    this_5_0_1_address0,
    this_5_0_1_ce0,
    this_5_0_1_we0,
    this_5_0_1_d0,
    this_5_0_1_q0,
    this_5_0_2_address0,
    this_5_0_2_ce0,
    this_5_0_2_we0,
    this_5_0_2_d0,
    this_5_0_2_q0,
    this_5_0_3_address0,
    this_5_0_3_ce0,
    this_5_0_3_we0,
    this_5_0_3_d0,
    this_5_0_3_q0,
    this_5_1_0_address0,
    this_5_1_0_ce0,
    this_5_1_0_we0,
    this_5_1_0_d0,
    this_5_1_0_q0,
    this_5_1_1_address0,
    this_5_1_1_ce0,
    this_5_1_1_we0,
    this_5_1_1_d0,
    this_5_1_1_q0,
    this_5_1_2_address0,
    this_5_1_2_ce0,
    this_5_1_2_we0,
    this_5_1_2_d0,
    this_5_1_2_q0,
    this_5_1_3_address0,
    this_5_1_3_ce0,
    this_5_1_3_we0,
    this_5_1_3_d0,
    this_5_1_3_q0,
    this_5_2_0_address0,
    this_5_2_0_ce0,
    this_5_2_0_we0,
    this_5_2_0_d0,
    this_5_2_0_q0,
    this_5_2_1_address0,
    this_5_2_1_ce0,
    this_5_2_1_we0,
    this_5_2_1_d0,
    this_5_2_1_q0,
    this_5_2_2_address0,
    this_5_2_2_ce0,
    this_5_2_2_we0,
    this_5_2_2_d0,
    this_5_2_2_q0,
    this_5_2_3_address0,
    this_5_2_3_ce0,
    this_5_2_3_we0,
    this_5_2_3_d0,
    this_5_2_3_q0,
    this_5_3_0_address0,
    this_5_3_0_ce0,
    this_5_3_0_we0,
    this_5_3_0_d0,
    this_5_3_0_q0,
    this_5_3_1_address0,
    this_5_3_1_ce0,
    this_5_3_1_we0,
    this_5_3_1_d0,
    this_5_3_1_q0,
    this_5_3_2_address0,
    this_5_3_2_ce0,
    this_5_3_2_we0,
    this_5_3_2_d0,
    this_5_3_2_q0,
    this_5_3_3_address0,
    this_5_3_3_ce0,
    this_5_3_3_we0,
    this_5_3_3_d0,
    this_5_3_3_q0,
    this_6_0_0_address0,
    this_6_0_0_ce0,
    this_6_0_0_we0,
    this_6_0_0_d0,
    this_6_0_0_q0,
    this_6_0_1_address0,
    this_6_0_1_ce0,
    this_6_0_1_we0,
    this_6_0_1_d0,
    this_6_0_1_q0,
    this_6_0_2_address0,
    this_6_0_2_ce0,
    this_6_0_2_we0,
    this_6_0_2_d0,
    this_6_0_2_q0,
    this_6_0_3_address0,
    this_6_0_3_ce0,
    this_6_0_3_we0,
    this_6_0_3_d0,
    this_6_0_3_q0,
    this_6_1_0_address0,
    this_6_1_0_ce0,
    this_6_1_0_we0,
    this_6_1_0_d0,
    this_6_1_0_q0,
    this_6_1_1_address0,
    this_6_1_1_ce0,
    this_6_1_1_we0,
    this_6_1_1_d0,
    this_6_1_1_q0,
    this_6_1_2_address0,
    this_6_1_2_ce0,
    this_6_1_2_we0,
    this_6_1_2_d0,
    this_6_1_2_q0,
    this_6_1_3_address0,
    this_6_1_3_ce0,
    this_6_1_3_we0,
    this_6_1_3_d0,
    this_6_1_3_q0,
    this_6_2_0_address0,
    this_6_2_0_ce0,
    this_6_2_0_we0,
    this_6_2_0_d0,
    this_6_2_0_q0,
    this_6_2_1_address0,
    this_6_2_1_ce0,
    this_6_2_1_we0,
    this_6_2_1_d0,
    this_6_2_1_q0,
    this_6_2_2_address0,
    this_6_2_2_ce0,
    this_6_2_2_we0,
    this_6_2_2_d0,
    this_6_2_2_q0,
    this_6_2_3_address0,
    this_6_2_3_ce0,
    this_6_2_3_we0,
    this_6_2_3_d0,
    this_6_2_3_q0,
    this_6_3_0_address0,
    this_6_3_0_ce0,
    this_6_3_0_we0,
    this_6_3_0_d0,
    this_6_3_0_q0,
    this_6_3_1_address0,
    this_6_3_1_ce0,
    this_6_3_1_we0,
    this_6_3_1_d0,
    this_6_3_1_q0,
    this_6_3_2_address0,
    this_6_3_2_ce0,
    this_6_3_2_we0,
    this_6_3_2_d0,
    this_6_3_2_q0,
    this_6_3_3_address0,
    this_6_3_3_ce0,
    this_6_3_3_we0,
    this_6_3_3_d0,
    this_6_3_3_q0,
    this_7_address0,
    this_7_ce0,
    this_7_we0,
    this_7_d0,
    this_7_q0,
    p_read,
    p_read1,
    p_read2,
    p_read3,
    p_read4,
    p_read5,
    p_read6,
    p_read7,
    p_read8,
    p_read9,
    p_read10,
    p_read11,
    p_read12,
    p_read13,
    p_read14,
    p_read15,
    p_read16,
    p_read17,
    p_read18,
    p_read19,
    p_read20,
    p_read21,
    p_read22,
    p_read23,
    p_read24,
    p_read25,
    p_read26,
    p_read27,
    p_read28,
    p_read29,
    p_read30,
    p_read31,
    p_read32,
    p_read33,
    p_read34,
    p_read35,
    p_read36,
    p_read37,
    p_read38,
    p_read39,
    p_read40,
    p_read41,
    p_read42,
    p_read43,
    p_read44,
    p_read45,
    p_read46,
    p_read47,
    p_read48,
    p_read49,
    p_read50,
    p_read51,
    p_read52,
    p_read53,
    p_read54,
    p_read55,
    p_read56,
    p_read57,
    p_read58,
    p_read59,
    p_read60,
    p_read61,
    p_read62,
    p_read63,
    this_15_address0,
    this_15_ce0,
    this_15_we0,
    this_15_d0,
    this_15_q0,
    this_15_address1,
    this_15_ce1,
    this_15_we1,
    this_15_d1,
    this_15_q1,
    this_16_address0,
    this_16_ce0,
    this_16_we0,
    this_16_d0,
    this_16_q0,
    this_16_address1,
    this_16_ce1,
    this_16_q1,
    l_TColl_0_0_0_constprop_i,
    l_TColl_0_0_0_constprop_o,
    l_TColl_0_0_0_constprop_o_ap_vld,
    l_TColl_0_0_1_constprop_i,
    l_TColl_0_0_1_constprop_o,
    l_TColl_0_0_1_constprop_o_ap_vld,
    l_TColl_0_0_2_constprop_i,
    l_TColl_0_0_2_constprop_o,
    l_TColl_0_0_2_constprop_o_ap_vld,
    l_TColl_0_0_3_constprop_i,
    l_TColl_0_0_3_constprop_o,
    l_TColl_0_0_3_constprop_o_ap_vld,
    l_TColl_1_0_0_constprop_i,
    l_TColl_1_0_0_constprop_o,
    l_TColl_1_0_0_constprop_o_ap_vld,
    l_TColl_1_0_1_constprop_i,
    l_TColl_1_0_1_constprop_o,
    l_TColl_1_0_1_constprop_o_ap_vld,
    l_TColl_1_0_2_constprop_i,
    l_TColl_1_0_2_constprop_o,
    l_TColl_1_0_2_constprop_o_ap_vld,
    l_TColl_1_0_3_constprop_i,
    l_TColl_1_0_3_constprop_o,
    l_TColl_1_0_3_constprop_o_ap_vld,
    l_TColl_2_0_0_constprop_i,
    l_TColl_2_0_0_constprop_o,
    l_TColl_2_0_0_constprop_o_ap_vld,
    l_TColl_2_0_1_constprop_i,
    l_TColl_2_0_1_constprop_o,
    l_TColl_2_0_1_constprop_o_ap_vld,
    l_TColl_2_0_2_constprop_i,
    l_TColl_2_0_2_constprop_o,
    l_TColl_2_0_2_constprop_o_ap_vld,
    l_TColl_2_0_3_constprop_i,
    l_TColl_2_0_3_constprop_o,
    l_TColl_2_0_3_constprop_o_ap_vld,
    l_TColl_0_1_0_constprop_i,
    l_TColl_0_1_0_constprop_o,
    l_TColl_0_1_0_constprop_o_ap_vld,
    l_TColl_0_1_1_constprop_i,
    l_TColl_0_1_1_constprop_o,
    l_TColl_0_1_1_constprop_o_ap_vld,
    l_TColl_0_1_2_constprop_i,
    l_TColl_0_1_2_constprop_o,
    l_TColl_0_1_2_constprop_o_ap_vld,
    l_TColl_0_1_3_constprop_i,
    l_TColl_0_1_3_constprop_o,
    l_TColl_0_1_3_constprop_o_ap_vld,
    l_TColl_1_1_0_constprop_i,
    l_TColl_1_1_0_constprop_o,
    l_TColl_1_1_0_constprop_o_ap_vld,
    l_TColl_1_1_1_constprop_i,
    l_TColl_1_1_1_constprop_o,
    l_TColl_1_1_1_constprop_o_ap_vld,
    l_TColl_1_1_2_constprop_i,
    l_TColl_1_1_2_constprop_o,
    l_TColl_1_1_2_constprop_o_ap_vld,
    l_TColl_1_1_3_constprop_i,
    l_TColl_1_1_3_constprop_o,
    l_TColl_1_1_3_constprop_o_ap_vld,
    l_TColl_2_1_0_constprop_i,
    l_TColl_2_1_0_constprop_o,
    l_TColl_2_1_0_constprop_o_ap_vld,
    l_TColl_2_1_1_constprop_i,
    l_TColl_2_1_1_constprop_o,
    l_TColl_2_1_1_constprop_o_ap_vld,
    l_TColl_2_1_2_constprop_i,
    l_TColl_2_1_2_constprop_o,
    l_TColl_2_1_2_constprop_o_ap_vld,
    l_TColl_2_1_3_constprop_i,
    l_TColl_2_1_3_constprop_o,
    l_TColl_2_1_3_constprop_o_ap_vld,
    l_TColl_0_2_0_constprop_i,
    l_TColl_0_2_0_constprop_o,
    l_TColl_0_2_0_constprop_o_ap_vld,
    l_TColl_0_2_1_constprop_i,
    l_TColl_0_2_1_constprop_o,
    l_TColl_0_2_1_constprop_o_ap_vld,
    l_TColl_0_2_2_constprop_i,
    l_TColl_0_2_2_constprop_o,
    l_TColl_0_2_2_constprop_o_ap_vld,
    l_TColl_0_2_3_constprop_i,
    l_TColl_0_2_3_constprop_o,
    l_TColl_0_2_3_constprop_o_ap_vld,
    l_TColl_1_2_0_constprop_i,
    l_TColl_1_2_0_constprop_o,
    l_TColl_1_2_0_constprop_o_ap_vld,
    l_TColl_1_2_1_constprop_i,
    l_TColl_1_2_1_constprop_o,
    l_TColl_1_2_1_constprop_o_ap_vld,
    l_TColl_1_2_2_constprop_i,
    l_TColl_1_2_2_constprop_o,
    l_TColl_1_2_2_constprop_o_ap_vld,
    l_TColl_1_2_3_constprop_i,
    l_TColl_1_2_3_constprop_o,
    l_TColl_1_2_3_constprop_o_ap_vld,
    l_TColl_2_2_0_constprop_i,
    l_TColl_2_2_0_constprop_o,
    l_TColl_2_2_0_constprop_o_ap_vld,
    l_TColl_2_2_1_constprop_i,
    l_TColl_2_2_1_constprop_o,
    l_TColl_2_2_1_constprop_o_ap_vld,
    l_TColl_2_2_2_constprop_i,
    l_TColl_2_2_2_constprop_o,
    l_TColl_2_2_2_constprop_o_ap_vld,
    l_TColl_2_2_3_constprop_i,
    l_TColl_2_2_3_constprop_o,
    l_TColl_2_2_3_constprop_o_ap_vld,
    l_TColl_0_3_0_constprop_i,
    l_TColl_0_3_0_constprop_o,
    l_TColl_0_3_0_constprop_o_ap_vld,
    l_TColl_0_3_1_constprop_i,
    l_TColl_0_3_1_constprop_o,
    l_TColl_0_3_1_constprop_o_ap_vld,
    l_TColl_0_3_2_constprop_i,
    l_TColl_0_3_2_constprop_o,
    l_TColl_0_3_2_constprop_o_ap_vld,
    l_TColl_0_3_3_constprop_i,
    l_TColl_0_3_3_constprop_o,
    l_TColl_0_3_3_constprop_o_ap_vld,
    l_TColl_1_3_0_constprop_i,
    l_TColl_1_3_0_constprop_o,
    l_TColl_1_3_0_constprop_o_ap_vld,
    l_TColl_1_3_1_constprop_i,
    l_TColl_1_3_1_constprop_o,
    l_TColl_1_3_1_constprop_o_ap_vld,
    l_TColl_1_3_2_constprop_i,
    l_TColl_1_3_2_constprop_o,
    l_TColl_1_3_2_constprop_o_ap_vld,
    l_TColl_1_3_3_constprop_i,
    l_TColl_1_3_3_constprop_o,
    l_TColl_1_3_3_constprop_o_ap_vld,
    l_TColl_2_3_0_constprop_i,
    l_TColl_2_3_0_constprop_o,
    l_TColl_2_3_0_constprop_o_ap_vld,
    l_TColl_2_3_1_constprop_i,
    l_TColl_2_3_1_constprop_o,
    l_TColl_2_3_1_constprop_o_ap_vld,
    l_TColl_2_3_2_constprop_i,
    l_TColl_2_3_2_constprop_o,
    l_TColl_2_3_2_constprop_o_ap_vld,
    l_TColl_2_3_3_constprop_i,
    l_TColl_2_3_3_constprop_o,
    l_TColl_2_3_3_constprop_o_ap_vld,
    grp_fu_2427_p_din0,
    grp_fu_2427_p_din1,
    grp_fu_2427_p_opcode,
    grp_fu_2427_p_dout0,
    grp_fu_2427_p_ce,
    grp_fu_2403_p_din0,
    grp_fu_2403_p_din1,
    grp_fu_2403_p_opcode,
    grp_fu_2403_p_dout0,
    grp_fu_2403_p_ce,
    grp_fu_2431_p_din0,
    grp_fu_2431_p_din1,
    grp_fu_2431_p_dout0,
    grp_fu_2431_p_ce,
    grp_fu_2407_p_din0,
    grp_fu_2407_p_din1,
    grp_fu_2407_p_opcode,
    grp_fu_2407_p_dout0,
    grp_fu_2407_p_ce,
    grp_fu_2411_p_din0,
    grp_fu_2411_p_din1,
    grp_fu_2411_p_opcode,
    grp_fu_2411_p_dout0,
    grp_fu_2411_p_ce,
    grp_fu_2415_p_din0,
    grp_fu_2415_p_din1,
    grp_fu_2415_p_opcode,
    grp_fu_2415_p_dout0,
    grp_fu_2415_p_ce,
    grp_fu_2419_p_din0,
    grp_fu_2419_p_din1,
    grp_fu_2419_p_opcode,
    grp_fu_2419_p_dout0,
    grp_fu_2419_p_ce,
    grp_fu_2423_p_din0,
    grp_fu_2423_p_din1,
    grp_fu_2423_p_opcode,
    grp_fu_2423_p_dout0,
    grp_fu_2423_p_ce,
    grp_fu_2435_p_din0,
    grp_fu_2435_p_din1,
    grp_fu_2435_p_dout0,
    grp_fu_2435_p_ce,
    grp_fu_2439_p_din0,
    grp_fu_2439_p_din1,
    grp_fu_2439_p_dout0,
    grp_fu_2439_p_ce,
    grp_fu_2443_p_din0,
    grp_fu_2443_p_din1,
    grp_fu_2443_p_dout0,
    grp_fu_2443_p_ce
);

    parameter ap_ST_fsm_state1 = 338'd1;
    parameter ap_ST_fsm_state2 = 338'd2;
    parameter ap_ST_fsm_state3 = 338'd4;
    parameter ap_ST_fsm_state4 = 338'd8;
    parameter ap_ST_fsm_state5 = 338'd16;
    parameter ap_ST_fsm_state6 = 338'd32;
    parameter ap_ST_fsm_state7 = 338'd64;
    parameter ap_ST_fsm_state8 = 338'd128;
    parameter ap_ST_fsm_state9 = 338'd256;
    parameter ap_ST_fsm_state10 = 338'd512;
    parameter ap_ST_fsm_state11 = 338'd1024;
    parameter ap_ST_fsm_state12 = 338'd2048;
    parameter ap_ST_fsm_state13 = 338'd4096;
    parameter ap_ST_fsm_state14 = 338'd8192;
    parameter ap_ST_fsm_state15 = 338'd16384;
    parameter ap_ST_fsm_state16 = 338'd32768;
    parameter ap_ST_fsm_state17 = 338'd65536;
    parameter ap_ST_fsm_state18 = 338'd131072;
    parameter ap_ST_fsm_state19 = 338'd262144;
    parameter ap_ST_fsm_state20 = 338'd524288;
    parameter ap_ST_fsm_state21 = 338'd1048576;
    parameter ap_ST_fsm_state22 = 338'd2097152;
    parameter ap_ST_fsm_state23 = 338'd4194304;
    parameter ap_ST_fsm_state24 = 338'd8388608;
    parameter ap_ST_fsm_state25 = 338'd16777216;
    parameter ap_ST_fsm_state26 = 338'd33554432;
    parameter ap_ST_fsm_state27 = 338'd67108864;
    parameter ap_ST_fsm_state28 = 338'd134217728;
    parameter ap_ST_fsm_state29 = 338'd268435456;
    parameter ap_ST_fsm_state30 = 338'd536870912;
    parameter ap_ST_fsm_state31 = 338'd1073741824;
    parameter ap_ST_fsm_state32 = 338'd2147483648;
    parameter ap_ST_fsm_state33 = 338'd4294967296;
    parameter ap_ST_fsm_state34 = 338'd8589934592;
    parameter ap_ST_fsm_state35 = 338'd17179869184;
    parameter ap_ST_fsm_state36 = 338'd34359738368;
    parameter ap_ST_fsm_state37 = 338'd68719476736;
    parameter ap_ST_fsm_state38 = 338'd137438953472;
    parameter ap_ST_fsm_state39 = 338'd274877906944;
    parameter ap_ST_fsm_state40 = 338'd549755813888;
    parameter ap_ST_fsm_state41 = 338'd1099511627776;
    parameter ap_ST_fsm_state42 = 338'd2199023255552;
    parameter ap_ST_fsm_state43 = 338'd4398046511104;
    parameter ap_ST_fsm_state44 = 338'd8796093022208;
    parameter ap_ST_fsm_state45 = 338'd17592186044416;
    parameter ap_ST_fsm_state46 = 338'd35184372088832;
    parameter ap_ST_fsm_state47 = 338'd70368744177664;
    parameter ap_ST_fsm_state48 = 338'd140737488355328;
    parameter ap_ST_fsm_state49 = 338'd281474976710656;
    parameter ap_ST_fsm_state50 = 338'd562949953421312;
    parameter ap_ST_fsm_state51 = 338'd1125899906842624;
    parameter ap_ST_fsm_state52 = 338'd2251799813685248;
    parameter ap_ST_fsm_state53 = 338'd4503599627370496;
    parameter ap_ST_fsm_state54 = 338'd9007199254740992;
    parameter ap_ST_fsm_state55 = 338'd18014398509481984;
    parameter ap_ST_fsm_state56 = 338'd36028797018963968;
    parameter ap_ST_fsm_state57 = 338'd72057594037927936;
    parameter ap_ST_fsm_state58 = 338'd144115188075855872;
    parameter ap_ST_fsm_state59 = 338'd288230376151711744;
    parameter ap_ST_fsm_state60 = 338'd576460752303423488;
    parameter ap_ST_fsm_state61 = 338'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 338'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 338'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 338'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 338'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 338'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 338'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 338'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 338'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 338'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 338'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 338'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 338'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 338'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 338'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 338'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 338'd75557863725914323419136;
    parameter ap_ST_fsm_state78 = 338'd151115727451828646838272;
    parameter ap_ST_fsm_state79 = 338'd302231454903657293676544;
    parameter ap_ST_fsm_state80 = 338'd604462909807314587353088;
    parameter ap_ST_fsm_state81 = 338'd1208925819614629174706176;
    parameter ap_ST_fsm_state82 = 338'd2417851639229258349412352;
    parameter ap_ST_fsm_state83 = 338'd4835703278458516698824704;
    parameter ap_ST_fsm_state84 = 338'd9671406556917033397649408;
    parameter ap_ST_fsm_state85 = 338'd19342813113834066795298816;
    parameter ap_ST_fsm_state86 = 338'd38685626227668133590597632;
    parameter ap_ST_fsm_state87 = 338'd77371252455336267181195264;
    parameter ap_ST_fsm_state88 = 338'd154742504910672534362390528;
    parameter ap_ST_fsm_state89 = 338'd309485009821345068724781056;
    parameter ap_ST_fsm_state90 = 338'd618970019642690137449562112;
    parameter ap_ST_fsm_state91 = 338'd1237940039285380274899124224;
    parameter ap_ST_fsm_state92 = 338'd2475880078570760549798248448;
    parameter ap_ST_fsm_state93 = 338'd4951760157141521099596496896;
    parameter ap_ST_fsm_state94 = 338'd9903520314283042199192993792;
    parameter ap_ST_fsm_state95 = 338'd19807040628566084398385987584;
    parameter ap_ST_fsm_state96 = 338'd39614081257132168796771975168;
    parameter ap_ST_fsm_state97 = 338'd79228162514264337593543950336;
    parameter ap_ST_fsm_state98 = 338'd158456325028528675187087900672;
    parameter ap_ST_fsm_state99 = 338'd316912650057057350374175801344;
    parameter ap_ST_fsm_state100 = 338'd633825300114114700748351602688;
    parameter ap_ST_fsm_state101 = 338'd1267650600228229401496703205376;
    parameter ap_ST_fsm_state102 = 338'd2535301200456458802993406410752;
    parameter ap_ST_fsm_state103 = 338'd5070602400912917605986812821504;
    parameter ap_ST_fsm_state104 = 338'd10141204801825835211973625643008;
    parameter ap_ST_fsm_state105 = 338'd20282409603651670423947251286016;
    parameter ap_ST_fsm_state106 = 338'd40564819207303340847894502572032;
    parameter ap_ST_fsm_state107 = 338'd81129638414606681695789005144064;
    parameter ap_ST_fsm_state108 = 338'd162259276829213363391578010288128;
    parameter ap_ST_fsm_state109 = 338'd324518553658426726783156020576256;
    parameter ap_ST_fsm_state110 = 338'd649037107316853453566312041152512;
    parameter ap_ST_fsm_state111 = 338'd1298074214633706907132624082305024;
    parameter ap_ST_fsm_state112 = 338'd2596148429267413814265248164610048;
    parameter ap_ST_fsm_state113 = 338'd5192296858534827628530496329220096;
    parameter ap_ST_fsm_state114 = 338'd10384593717069655257060992658440192;
    parameter ap_ST_fsm_state115 = 338'd20769187434139310514121985316880384;
    parameter ap_ST_fsm_state116 = 338'd41538374868278621028243970633760768;
    parameter ap_ST_fsm_state117 = 338'd83076749736557242056487941267521536;
    parameter ap_ST_fsm_state118 = 338'd166153499473114484112975882535043072;
    parameter ap_ST_fsm_state119 = 338'd332306998946228968225951765070086144;
    parameter ap_ST_fsm_state120 = 338'd664613997892457936451903530140172288;
    parameter ap_ST_fsm_state121 = 338'd1329227995784915872903807060280344576;
    parameter ap_ST_fsm_state122 = 338'd2658455991569831745807614120560689152;
    parameter ap_ST_fsm_state123 = 338'd5316911983139663491615228241121378304;
    parameter ap_ST_fsm_state124 = 338'd10633823966279326983230456482242756608;
    parameter ap_ST_fsm_state125 = 338'd21267647932558653966460912964485513216;
    parameter ap_ST_fsm_state126 = 338'd42535295865117307932921825928971026432;
    parameter ap_ST_fsm_state127 = 338'd85070591730234615865843651857942052864;
    parameter ap_ST_fsm_state128 = 338'd170141183460469231731687303715884105728;
    parameter ap_ST_fsm_state129 = 338'd340282366920938463463374607431768211456;
    parameter ap_ST_fsm_state130 = 338'd680564733841876926926749214863536422912;
    parameter ap_ST_fsm_state131 = 338'd1361129467683753853853498429727072845824;
    parameter ap_ST_fsm_state132 = 338'd2722258935367507707706996859454145691648;
    parameter ap_ST_fsm_state133 = 338'd5444517870735015415413993718908291383296;
    parameter ap_ST_fsm_state134 = 338'd10889035741470030830827987437816582766592;
    parameter ap_ST_fsm_state135 = 338'd21778071482940061661655974875633165533184;
    parameter ap_ST_fsm_state136 = 338'd43556142965880123323311949751266331066368;
    parameter ap_ST_fsm_state137 = 338'd87112285931760246646623899502532662132736;
    parameter ap_ST_fsm_state138 = 338'd174224571863520493293247799005065324265472;
    parameter ap_ST_fsm_state139 = 338'd348449143727040986586495598010130648530944;
    parameter ap_ST_fsm_state140 = 338'd696898287454081973172991196020261297061888;
    parameter ap_ST_fsm_state141 = 338'd1393796574908163946345982392040522594123776;
    parameter ap_ST_fsm_state142 = 338'd2787593149816327892691964784081045188247552;
    parameter ap_ST_fsm_state143 = 338'd5575186299632655785383929568162090376495104;
    parameter ap_ST_fsm_state144 = 338'd11150372599265311570767859136324180752990208;
    parameter ap_ST_fsm_state145 = 338'd22300745198530623141535718272648361505980416;
    parameter ap_ST_fsm_state146 = 338'd44601490397061246283071436545296723011960832;
    parameter ap_ST_fsm_state147 = 338'd89202980794122492566142873090593446023921664;
    parameter ap_ST_fsm_state148 = 338'd178405961588244985132285746181186892047843328;
    parameter ap_ST_fsm_state149 = 338'd356811923176489970264571492362373784095686656;
    parameter ap_ST_fsm_state150 = 338'd713623846352979940529142984724747568191373312;
    parameter ap_ST_fsm_state151 = 338'd1427247692705959881058285969449495136382746624;
    parameter ap_ST_fsm_state152 = 338'd2854495385411919762116571938898990272765493248;
    parameter ap_ST_fsm_state153 = 338'd5708990770823839524233143877797980545530986496;
    parameter ap_ST_fsm_state154 = 338'd11417981541647679048466287755595961091061972992;
    parameter ap_ST_fsm_state155 = 338'd22835963083295358096932575511191922182123945984;
    parameter ap_ST_fsm_state156 = 338'd45671926166590716193865151022383844364247891968;
    parameter ap_ST_fsm_state157 = 338'd91343852333181432387730302044767688728495783936;
    parameter ap_ST_fsm_state158 = 338'd182687704666362864775460604089535377456991567872;
    parameter ap_ST_fsm_state159 = 338'd365375409332725729550921208179070754913983135744;
    parameter ap_ST_fsm_state160 = 338'd730750818665451459101842416358141509827966271488;
    parameter ap_ST_fsm_state161 = 338'd1461501637330902918203684832716283019655932542976;
    parameter ap_ST_fsm_state162 = 338'd2923003274661805836407369665432566039311865085952;
    parameter ap_ST_fsm_state163 = 338'd5846006549323611672814739330865132078623730171904;
    parameter ap_ST_fsm_state164 = 338'd11692013098647223345629478661730264157247460343808;
    parameter ap_ST_fsm_state165 = 338'd23384026197294446691258957323460528314494920687616;
    parameter ap_ST_fsm_state166 = 338'd46768052394588893382517914646921056628989841375232;
    parameter ap_ST_fsm_state167 = 338'd93536104789177786765035829293842113257979682750464;
    parameter ap_ST_fsm_state168 = 338'd187072209578355573530071658587684226515959365500928;
    parameter ap_ST_fsm_state169 = 338'd374144419156711147060143317175368453031918731001856;
    parameter ap_ST_fsm_state170 = 338'd748288838313422294120286634350736906063837462003712;
    parameter ap_ST_fsm_state171 = 338'd1496577676626844588240573268701473812127674924007424;
    parameter ap_ST_fsm_state172 = 338'd2993155353253689176481146537402947624255349848014848;
    parameter ap_ST_fsm_state173 = 338'd5986310706507378352962293074805895248510699696029696;
    parameter ap_ST_fsm_state174 = 338'd11972621413014756705924586149611790497021399392059392;
    parameter ap_ST_fsm_state175 = 338'd23945242826029513411849172299223580994042798784118784;
    parameter ap_ST_fsm_state176 = 338'd47890485652059026823698344598447161988085597568237568;
    parameter ap_ST_fsm_state177 = 338'd95780971304118053647396689196894323976171195136475136;
    parameter ap_ST_fsm_state178 = 338'd191561942608236107294793378393788647952342390272950272;
    parameter ap_ST_fsm_state179 = 338'd383123885216472214589586756787577295904684780545900544;
    parameter ap_ST_fsm_state180 = 338'd766247770432944429179173513575154591809369561091801088;
    parameter ap_ST_fsm_state181 = 338'd1532495540865888858358347027150309183618739122183602176;
    parameter ap_ST_fsm_state182 = 338'd3064991081731777716716694054300618367237478244367204352;
    parameter ap_ST_fsm_state183 = 338'd6129982163463555433433388108601236734474956488734408704;
    parameter ap_ST_fsm_state184 = 338'd12259964326927110866866776217202473468949912977468817408;
    parameter ap_ST_fsm_state185 = 338'd24519928653854221733733552434404946937899825954937634816;
    parameter ap_ST_fsm_state186 = 338'd49039857307708443467467104868809893875799651909875269632;
    parameter ap_ST_fsm_state187 = 338'd98079714615416886934934209737619787751599303819750539264;
    parameter ap_ST_fsm_state188 = 338'd196159429230833773869868419475239575503198607639501078528;
    parameter ap_ST_fsm_state189 = 338'd392318858461667547739736838950479151006397215279002157056;
    parameter ap_ST_fsm_state190 = 338'd784637716923335095479473677900958302012794430558004314112;
    parameter ap_ST_fsm_state191 = 338'd1569275433846670190958947355801916604025588861116008628224;
    parameter ap_ST_fsm_state192 = 338'd3138550867693340381917894711603833208051177722232017256448;
    parameter ap_ST_fsm_state193 = 338'd6277101735386680763835789423207666416102355444464034512896;
    parameter ap_ST_fsm_state194 = 338'd12554203470773361527671578846415332832204710888928069025792;
    parameter ap_ST_fsm_state195 = 338'd25108406941546723055343157692830665664409421777856138051584;
    parameter ap_ST_fsm_state196 = 338'd50216813883093446110686315385661331328818843555712276103168;
    parameter    ap_ST_fsm_state197 = 338'd100433627766186892221372630771322662657637687111424552206336;
    parameter    ap_ST_fsm_state198 = 338'd200867255532373784442745261542645325315275374222849104412672;
    parameter    ap_ST_fsm_state199 = 338'd401734511064747568885490523085290650630550748445698208825344;
    parameter    ap_ST_fsm_state200 = 338'd803469022129495137770981046170581301261101496891396417650688;
    parameter    ap_ST_fsm_state201 = 338'd1606938044258990275541962092341162602522202993782792835301376;
    parameter    ap_ST_fsm_state202 = 338'd3213876088517980551083924184682325205044405987565585670602752;
    parameter    ap_ST_fsm_state203 = 338'd6427752177035961102167848369364650410088811975131171341205504;
    parameter    ap_ST_fsm_state204 = 338'd12855504354071922204335696738729300820177623950262342682411008;
    parameter    ap_ST_fsm_state205 = 338'd25711008708143844408671393477458601640355247900524685364822016;
    parameter    ap_ST_fsm_state206 = 338'd51422017416287688817342786954917203280710495801049370729644032;
    parameter    ap_ST_fsm_state207 = 338'd102844034832575377634685573909834406561420991602098741459288064;
    parameter    ap_ST_fsm_state208 = 338'd205688069665150755269371147819668813122841983204197482918576128;
    parameter    ap_ST_fsm_state209 = 338'd411376139330301510538742295639337626245683966408394965837152256;
    parameter    ap_ST_fsm_state210 = 338'd822752278660603021077484591278675252491367932816789931674304512;
    parameter    ap_ST_fsm_state211 = 338'd1645504557321206042154969182557350504982735865633579863348609024;
    parameter    ap_ST_fsm_state212 = 338'd3291009114642412084309938365114701009965471731267159726697218048;
    parameter    ap_ST_fsm_state213 = 338'd6582018229284824168619876730229402019930943462534319453394436096;
    parameter    ap_ST_fsm_state214 = 338'd13164036458569648337239753460458804039861886925068638906788872192;
    parameter    ap_ST_fsm_state215 = 338'd26328072917139296674479506920917608079723773850137277813577744384;
    parameter    ap_ST_fsm_state216 = 338'd52656145834278593348959013841835216159447547700274555627155488768;
    parameter    ap_ST_fsm_state217 = 338'd105312291668557186697918027683670432318895095400549111254310977536;
    parameter    ap_ST_fsm_state218 = 338'd210624583337114373395836055367340864637790190801098222508621955072;
    parameter    ap_ST_fsm_state219 = 338'd421249166674228746791672110734681729275580381602196445017243910144;
    parameter    ap_ST_fsm_state220 = 338'd842498333348457493583344221469363458551160763204392890034487820288;
    parameter    ap_ST_fsm_state221 = 338'd1684996666696914987166688442938726917102321526408785780068975640576;
    parameter    ap_ST_fsm_state222 = 338'd3369993333393829974333376885877453834204643052817571560137951281152;
    parameter    ap_ST_fsm_state223 = 338'd6739986666787659948666753771754907668409286105635143120275902562304;
    parameter    ap_ST_fsm_state224 = 338'd13479973333575319897333507543509815336818572211270286240551805124608;
    parameter    ap_ST_fsm_state225 = 338'd26959946667150639794667015087019630673637144422540572481103610249216;
    parameter    ap_ST_fsm_state226 = 338'd53919893334301279589334030174039261347274288845081144962207220498432;
    parameter    ap_ST_fsm_state227 = 338'd107839786668602559178668060348078522694548577690162289924414440996864;
    parameter    ap_ST_fsm_state228 = 338'd215679573337205118357336120696157045389097155380324579848828881993728;
    parameter    ap_ST_fsm_state229 = 338'd431359146674410236714672241392314090778194310760649159697657763987456;
    parameter    ap_ST_fsm_state230 = 338'd862718293348820473429344482784628181556388621521298319395315527974912;
    parameter    ap_ST_fsm_state231 = 338'd1725436586697640946858688965569256363112777243042596638790631055949824;
    parameter    ap_ST_fsm_state232 = 338'd3450873173395281893717377931138512726225554486085193277581262111899648;
    parameter    ap_ST_fsm_state233 = 338'd6901746346790563787434755862277025452451108972170386555162524223799296;
    parameter    ap_ST_fsm_state234 = 338'd13803492693581127574869511724554050904902217944340773110325048447598592;
    parameter    ap_ST_fsm_state235 = 338'd27606985387162255149739023449108101809804435888681546220650096895197184;
    parameter    ap_ST_fsm_state236 = 338'd55213970774324510299478046898216203619608871777363092441300193790394368;
    parameter    ap_ST_fsm_state237 = 338'd110427941548649020598956093796432407239217743554726184882600387580788736;
    parameter    ap_ST_fsm_state238 = 338'd220855883097298041197912187592864814478435487109452369765200775161577472;
    parameter    ap_ST_fsm_state239 = 338'd441711766194596082395824375185729628956870974218904739530401550323154944;
    parameter    ap_ST_fsm_state240 = 338'd883423532389192164791648750371459257913741948437809479060803100646309888;
    parameter    ap_ST_fsm_state241 = 338'd1766847064778384329583297500742918515827483896875618958121606201292619776;
    parameter    ap_ST_fsm_state242 = 338'd3533694129556768659166595001485837031654967793751237916243212402585239552;
    parameter    ap_ST_fsm_state243 = 338'd7067388259113537318333190002971674063309935587502475832486424805170479104;
    parameter    ap_ST_fsm_state244 = 338'd14134776518227074636666380005943348126619871175004951664972849610340958208;
    parameter    ap_ST_fsm_state245 = 338'd28269553036454149273332760011886696253239742350009903329945699220681916416;
    parameter    ap_ST_fsm_state246 = 338'd56539106072908298546665520023773392506479484700019806659891398441363832832;
    parameter    ap_ST_fsm_state247 = 338'd113078212145816597093331040047546785012958969400039613319782796882727665664;
    parameter    ap_ST_fsm_state248 = 338'd226156424291633194186662080095093570025917938800079226639565593765455331328;
    parameter    ap_ST_fsm_state249 = 338'd452312848583266388373324160190187140051835877600158453279131187530910662656;
    parameter    ap_ST_fsm_state250 = 338'd904625697166532776746648320380374280103671755200316906558262375061821325312;
    parameter    ap_ST_fsm_state251 = 338'd1809251394333065553493296640760748560207343510400633813116524750123642650624;
    parameter    ap_ST_fsm_state252 = 338'd3618502788666131106986593281521497120414687020801267626233049500247285301248;
    parameter    ap_ST_fsm_state253 = 338'd7237005577332262213973186563042994240829374041602535252466099000494570602496;
    parameter    ap_ST_fsm_state254 = 338'd14474011154664524427946373126085988481658748083205070504932198000989141204992;
    parameter    ap_ST_fsm_state255 = 338'd28948022309329048855892746252171976963317496166410141009864396001978282409984;
    parameter    ap_ST_fsm_state256 = 338'd57896044618658097711785492504343953926634992332820282019728792003956564819968;
    parameter    ap_ST_fsm_state257 = 338'd115792089237316195423570985008687907853269984665640564039457584007913129639936;
    parameter    ap_ST_fsm_state258 = 338'd231584178474632390847141970017375815706539969331281128078915168015826259279872;
    parameter    ap_ST_fsm_state259 = 338'd463168356949264781694283940034751631413079938662562256157830336031652518559744;
    parameter    ap_ST_fsm_state260 = 338'd926336713898529563388567880069503262826159877325124512315660672063305037119488;
    parameter    ap_ST_fsm_state261 = 338'd1852673427797059126777135760139006525652319754650249024631321344126610074238976;
    parameter    ap_ST_fsm_state262 = 338'd3705346855594118253554271520278013051304639509300498049262642688253220148477952;
    parameter    ap_ST_fsm_state263 = 338'd7410693711188236507108543040556026102609279018600996098525285376506440296955904;
    parameter    ap_ST_fsm_state264 = 338'd14821387422376473014217086081112052205218558037201992197050570753012880593911808;
    parameter    ap_ST_fsm_state265 = 338'd29642774844752946028434172162224104410437116074403984394101141506025761187823616;
    parameter    ap_ST_fsm_state266 = 338'd59285549689505892056868344324448208820874232148807968788202283012051522375647232;
    parameter    ap_ST_fsm_state267 = 338'd118571099379011784113736688648896417641748464297615937576404566024103044751294464;
    parameter    ap_ST_fsm_state268 = 338'd237142198758023568227473377297792835283496928595231875152809132048206089502588928;
    parameter    ap_ST_fsm_state269 = 338'd474284397516047136454946754595585670566993857190463750305618264096412179005177856;
    parameter    ap_ST_fsm_state270 = 338'd948568795032094272909893509191171341133987714380927500611236528192824358010355712;
    parameter    ap_ST_fsm_state271 = 338'd1897137590064188545819787018382342682267975428761855001222473056385648716020711424;
    parameter    ap_ST_fsm_state272 = 338'd3794275180128377091639574036764685364535950857523710002444946112771297432041422848;
    parameter    ap_ST_fsm_state273 = 338'd7588550360256754183279148073529370729071901715047420004889892225542594864082845696;
    parameter    ap_ST_fsm_state274 = 338'd15177100720513508366558296147058741458143803430094840009779784451085189728165691392;
    parameter    ap_ST_fsm_state275 = 338'd30354201441027016733116592294117482916287606860189680019559568902170379456331382784;
    parameter    ap_ST_fsm_state276 = 338'd60708402882054033466233184588234965832575213720379360039119137804340758912662765568;
    parameter    ap_ST_fsm_state277 = 338'd121416805764108066932466369176469931665150427440758720078238275608681517825325531136;
    parameter    ap_ST_fsm_state278 = 338'd242833611528216133864932738352939863330300854881517440156476551217363035650651062272;
    parameter    ap_ST_fsm_state279 = 338'd485667223056432267729865476705879726660601709763034880312953102434726071301302124544;
    parameter    ap_ST_fsm_state280 = 338'd971334446112864535459730953411759453321203419526069760625906204869452142602604249088;
    parameter    ap_ST_fsm_state281 = 338'd1942668892225729070919461906823518906642406839052139521251812409738904285205208498176;
    parameter    ap_ST_fsm_state282 = 338'd3885337784451458141838923813647037813284813678104279042503624819477808570410416996352;
    parameter    ap_ST_fsm_state283 = 338'd7770675568902916283677847627294075626569627356208558085007249638955617140820833992704;
    parameter    ap_ST_fsm_state284 = 338'd15541351137805832567355695254588151253139254712417116170014499277911234281641667985408;
    parameter    ap_ST_fsm_state285 = 338'd31082702275611665134711390509176302506278509424834232340028998555822468563283335970816;
    parameter    ap_ST_fsm_state286 = 338'd62165404551223330269422781018352605012557018849668464680057997111644937126566671941632;
    parameter    ap_ST_fsm_state287 = 338'd124330809102446660538845562036705210025114037699336929360115994223289874253133343883264;
    parameter    ap_ST_fsm_state288 = 338'd248661618204893321077691124073410420050228075398673858720231988446579748506266687766528;
    parameter    ap_ST_fsm_state289 = 338'd497323236409786642155382248146820840100456150797347717440463976893159497012533375533056;
    parameter    ap_ST_fsm_state290 = 338'd994646472819573284310764496293641680200912301594695434880927953786318994025066751066112;
    parameter    ap_ST_fsm_state291 = 338'd1989292945639146568621528992587283360401824603189390869761855907572637988050133502132224;
    parameter    ap_ST_fsm_state292 = 338'd3978585891278293137243057985174566720803649206378781739523711815145275976100267004264448;
    parameter    ap_ST_fsm_state293 = 338'd7957171782556586274486115970349133441607298412757563479047423630290551952200534008528896;
    parameter    ap_ST_fsm_state294 = 338'd15914343565113172548972231940698266883214596825515126958094847260581103904401068017057792;
    parameter    ap_ST_fsm_state295 = 338'd31828687130226345097944463881396533766429193651030253916189694521162207808802136034115584;
    parameter    ap_ST_fsm_state296 = 338'd63657374260452690195888927762793067532858387302060507832379389042324415617604272068231168;
    parameter    ap_ST_fsm_state297 = 338'd127314748520905380391777855525586135065716774604121015664758778084648831235208544136462336;
    parameter    ap_ST_fsm_state298 = 338'd254629497041810760783555711051172270131433549208242031329517556169297662470417088272924672;
    parameter    ap_ST_fsm_state299 = 338'd509258994083621521567111422102344540262867098416484062659035112338595324940834176545849344;
    parameter    ap_ST_fsm_state300 = 338'd1018517988167243043134222844204689080525734196832968125318070224677190649881668353091698688;
    parameter    ap_ST_fsm_state301 = 338'd2037035976334486086268445688409378161051468393665936250636140449354381299763336706183397376;
    parameter    ap_ST_fsm_state302 = 338'd4074071952668972172536891376818756322102936787331872501272280898708762599526673412366794752;
    parameter    ap_ST_fsm_state303 = 338'd8148143905337944345073782753637512644205873574663745002544561797417525199053346824733589504;
    parameter    ap_ST_fsm_state304 = 338'd16296287810675888690147565507275025288411747149327490005089123594835050398106693649467179008;
    parameter    ap_ST_fsm_state305 = 338'd32592575621351777380295131014550050576823494298654980010178247189670100796213387298934358016;
    parameter    ap_ST_fsm_state306 = 338'd65185151242703554760590262029100101153646988597309960020356494379340201592426774597868716032;
    parameter    ap_ST_fsm_state307 = 338'd130370302485407109521180524058200202307293977194619920040712988758680403184853549195737432064;
    parameter    ap_ST_fsm_state308 = 338'd260740604970814219042361048116400404614587954389239840081425977517360806369707098391474864128;
    parameter    ap_ST_fsm_state309 = 338'd521481209941628438084722096232800809229175908778479680162851955034721612739414196782949728256;
    parameter    ap_ST_fsm_state310 = 338'd1042962419883256876169444192465601618458351817556959360325703910069443225478828393565899456512;
    parameter    ap_ST_fsm_state311 = 338'd2085924839766513752338888384931203236916703635113918720651407820138886450957656787131798913024;
    parameter    ap_ST_fsm_state312 = 338'd4171849679533027504677776769862406473833407270227837441302815640277772901915313574263597826048;
    parameter    ap_ST_fsm_state313 = 338'd8343699359066055009355553539724812947666814540455674882605631280555545803830627148527195652096;
    parameter    ap_ST_fsm_state314 = 338'd16687398718132110018711107079449625895333629080911349765211262561111091607661254297054391304192;
    parameter    ap_ST_fsm_state315 = 338'd33374797436264220037422214158899251790667258161822699530422525122222183215322508594108782608384;
    parameter    ap_ST_fsm_state316 = 338'd66749594872528440074844428317798503581334516323645399060845050244444366430645017188217565216768;
    parameter    ap_ST_fsm_state317 = 338'd133499189745056880149688856635597007162669032647290798121690100488888732861290034376435130433536;
    parameter    ap_ST_fsm_state318 = 338'd266998379490113760299377713271194014325338065294581596243380200977777465722580068752870260867072;
    parameter    ap_ST_fsm_state319 = 338'd533996758980227520598755426542388028650676130589163192486760401955554931445160137505740521734144;
    parameter    ap_ST_fsm_state320 = 338'd1067993517960455041197510853084776057301352261178326384973520803911109862890320275011481043468288;
    parameter    ap_ST_fsm_state321 = 338'd2135987035920910082395021706169552114602704522356652769947041607822219725780640550022962086936576;
    parameter    ap_ST_fsm_state322 = 338'd4271974071841820164790043412339104229205409044713305539894083215644439451561281100045924173873152;
    parameter    ap_ST_fsm_state323 = 338'd8543948143683640329580086824678208458410818089426611079788166431288878903122562200091848347746304;
    parameter    ap_ST_fsm_state324 = 338'd17087896287367280659160173649356416916821636178853222159576332862577757806245124400183696695492608;
    parameter    ap_ST_fsm_state325 = 338'd34175792574734561318320347298712833833643272357706444319152665725155515612490248800367393390985216;
    parameter    ap_ST_fsm_state326 = 338'd68351585149469122636640694597425667667286544715412888638305331450311031224980497600734786781970432;
    parameter    ap_ST_fsm_state327 = 338'd136703170298938245273281389194851335334573089430825777276610662900622062449960995201469573563940864;
    parameter    ap_ST_fsm_state328 = 338'd273406340597876490546562778389702670669146178861651554553221325801244124899921990402939147127881728;
    parameter    ap_ST_fsm_state329 = 338'd546812681195752981093125556779405341338292357723303109106442651602488249799843980805878294255763456;
    parameter    ap_ST_fsm_state330 = 338'd1093625362391505962186251113558810682676584715446606218212885303204976499599687961611756588511526912;
    parameter    ap_ST_fsm_state331 = 338'd2187250724783011924372502227117621365353169430893212436425770606409952999199375923223513177023053824;
    parameter    ap_ST_fsm_state332 = 338'd4374501449566023848745004454235242730706338861786424872851541212819905998398751846447026354046107648;
    parameter    ap_ST_fsm_state333 = 338'd8749002899132047697490008908470485461412677723572849745703082425639811996797503692894052708092215296;
    parameter    ap_ST_fsm_state334 = 338'd17498005798264095394980017816940970922825355447145699491406164851279623993595007385788105416184430592;
    parameter    ap_ST_fsm_state335 = 338'd34996011596528190789960035633881941845650710894291398982812329702559247987190014771576210832368861184;
    parameter    ap_ST_fsm_state336 = 338'd69992023193056381579920071267763883691301421788582797965624659405118495974380029543152421664737722368;
    parameter    ap_ST_fsm_state337 = 338'd139984046386112763159840142535527767382602843577165595931249318810236991948760059086304843329475444736;
    parameter    ap_ST_fsm_state338 = 338'd279968092772225526319680285071055534765205687154331191862498637620473983897520118172609686658950889472;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [2:0] this_0_0_0_0_address0;
    output this_0_0_0_0_ce0;
    input [63:0] this_0_0_0_0_q0;
    output [2:0] this_0_0_0_1_address0;
    output this_0_0_0_1_ce0;
    input [63:0] this_0_0_0_1_q0;
    output [2:0] this_0_0_0_2_address0;
    output this_0_0_0_2_ce0;
    input [63:0] this_0_0_0_2_q0;
    output [2:0] this_0_0_1_0_address0;
    output this_0_0_1_0_ce0;
    input [63:0] this_0_0_1_0_q0;
    output [2:0] this_0_0_1_1_address0;
    output this_0_0_1_1_ce0;
    input [63:0] this_0_0_1_1_q0;
    output [2:0] this_0_0_1_2_address0;
    output this_0_0_1_2_ce0;
    input [63:0] this_0_0_1_2_q0;
    output [2:0] this_0_0_2_0_address0;
    output this_0_0_2_0_ce0;
    input [63:0] this_0_0_2_0_q0;
    output [2:0] this_0_0_2_1_address0;
    output this_0_0_2_1_ce0;
    input [63:0] this_0_0_2_1_q0;
    output [2:0] this_0_0_2_2_address0;
    output this_0_0_2_2_ce0;
    input [63:0] this_0_0_2_2_q0;
    output [2:0] this_0_0_3_0_address0;
    output this_0_0_3_0_ce0;
    input [63:0] this_0_0_3_0_q0;
    output [2:0] this_0_0_3_1_address0;
    output this_0_0_3_1_ce0;
    input [63:0] this_0_0_3_1_q0;
    output [2:0] this_0_0_3_2_address0;
    output this_0_0_3_2_ce0;
    input [63:0] this_0_0_3_2_q0;
    output [2:0] this_0_0_4_0_address0;
    output this_0_0_4_0_ce0;
    input [63:0] this_0_0_4_0_q0;
    output [2:0] this_0_0_4_1_address0;
    output this_0_0_4_1_ce0;
    input [63:0] this_0_0_4_1_q0;
    output [2:0] this_0_0_4_2_address0;
    output this_0_0_4_2_ce0;
    input [63:0] this_0_0_4_2_q0;
    output [2:0] this_0_0_5_0_address0;
    output this_0_0_5_0_ce0;
    input [63:0] this_0_0_5_0_q0;
    output [2:0] this_0_0_5_1_address0;
    output this_0_0_5_1_ce0;
    input [63:0] this_0_0_5_1_q0;
    output [2:0] this_0_0_5_2_address0;
    output this_0_0_5_2_ce0;
    input [63:0] this_0_0_5_2_q0;
    output [2:0] this_0_0_6_0_address0;
    output this_0_0_6_0_ce0;
    input [63:0] this_0_0_6_0_q0;
    output [2:0] this_0_0_6_1_address0;
    output this_0_0_6_1_ce0;
    input [63:0] this_0_0_6_1_q0;
    output [2:0] this_0_0_6_2_address0;
    output this_0_0_6_2_ce0;
    input [63:0] this_0_0_6_2_q0;
    output [2:0] this_0_0_7_0_address0;
    output this_0_0_7_0_ce0;
    input [63:0] this_0_0_7_0_q0;
    output [2:0] this_0_0_7_1_address0;
    output this_0_0_7_1_ce0;
    input [63:0] this_0_0_7_1_q0;
    output [2:0] this_0_0_7_2_address0;
    output this_0_0_7_2_ce0;
    input [63:0] this_0_0_7_2_q0;
    output [2:0] this_0_0_8_0_address0;
    output this_0_0_8_0_ce0;
    input [63:0] this_0_0_8_0_q0;
    output [2:0] this_0_0_8_1_address0;
    output this_0_0_8_1_ce0;
    input [63:0] this_0_0_8_1_q0;
    output [2:0] this_0_0_8_2_address0;
    output this_0_0_8_2_ce0;
    input [63:0] this_0_0_8_2_q0;
    output [6:0] this_0_1_address0;
    output this_0_1_ce0;
    input [63:0] this_0_1_q0;
    output [6:0] this_0_1_address1;
    output this_0_1_ce1;
    input [63:0] this_0_1_q1;
    output [2:0] this_4_0_0_address0;
    output this_4_0_0_ce0;
    input [63:0] this_4_0_0_q0;
    output [2:0] this_4_0_1_address0;
    output this_4_0_1_ce0;
    input [63:0] this_4_0_1_q0;
    output [2:0] this_4_0_2_address0;
    output this_4_0_2_ce0;
    input [63:0] this_4_0_2_q0;
    output [2:0] this_4_0_3_address0;
    output this_4_0_3_ce0;
    input [63:0] this_4_0_3_q0;
    output [2:0] this_4_1_0_address0;
    output this_4_1_0_ce0;
    input [63:0] this_4_1_0_q0;
    output [2:0] this_4_1_1_address0;
    output this_4_1_1_ce0;
    input [63:0] this_4_1_1_q0;
    output [2:0] this_4_1_2_address0;
    output this_4_1_2_ce0;
    input [63:0] this_4_1_2_q0;
    output [2:0] this_4_1_3_address0;
    output this_4_1_3_ce0;
    input [63:0] this_4_1_3_q0;
    output [2:0] this_4_2_0_address0;
    output this_4_2_0_ce0;
    input [63:0] this_4_2_0_q0;
    output [2:0] this_4_2_1_address0;
    output this_4_2_1_ce0;
    input [63:0] this_4_2_1_q0;
    output [2:0] this_4_2_2_address0;
    output this_4_2_2_ce0;
    input [63:0] this_4_2_2_q0;
    output [2:0] this_4_2_3_address0;
    output this_4_2_3_ce0;
    input [63:0] this_4_2_3_q0;
    output [2:0] this_4_3_0_address0;
    output this_4_3_0_ce0;
    input [63:0] this_4_3_0_q0;
    output [2:0] this_4_3_1_address0;
    output this_4_3_1_ce0;
    input [63:0] this_4_3_1_q0;
    output [2:0] this_4_3_2_address0;
    output this_4_3_2_ce0;
    input [63:0] this_4_3_2_q0;
    output [2:0] this_4_3_3_address0;
    output this_4_3_3_ce0;
    input [63:0] this_4_3_3_q0;
    output [2:0] this_5_0_0_address0;
    output this_5_0_0_ce0;
    output this_5_0_0_we0;
    output [63:0] this_5_0_0_d0;
    input [63:0] this_5_0_0_q0;
    output [2:0] this_5_0_1_address0;
    output this_5_0_1_ce0;
    output this_5_0_1_we0;
    output [63:0] this_5_0_1_d0;
    input [63:0] this_5_0_1_q0;
    output [2:0] this_5_0_2_address0;
    output this_5_0_2_ce0;
    output this_5_0_2_we0;
    output [63:0] this_5_0_2_d0;
    input [63:0] this_5_0_2_q0;
    output [2:0] this_5_0_3_address0;
    output this_5_0_3_ce0;
    output this_5_0_3_we0;
    output [63:0] this_5_0_3_d0;
    input [63:0] this_5_0_3_q0;
    output [2:0] this_5_1_0_address0;
    output this_5_1_0_ce0;
    output this_5_1_0_we0;
    output [63:0] this_5_1_0_d0;
    input [63:0] this_5_1_0_q0;
    output [2:0] this_5_1_1_address0;
    output this_5_1_1_ce0;
    output this_5_1_1_we0;
    output [63:0] this_5_1_1_d0;
    input [63:0] this_5_1_1_q0;
    output [2:0] this_5_1_2_address0;
    output this_5_1_2_ce0;
    output this_5_1_2_we0;
    output [63:0] this_5_1_2_d0;
    input [63:0] this_5_1_2_q0;
    output [2:0] this_5_1_3_address0;
    output this_5_1_3_ce0;
    output this_5_1_3_we0;
    output [63:0] this_5_1_3_d0;
    input [63:0] this_5_1_3_q0;
    output [2:0] this_5_2_0_address0;
    output this_5_2_0_ce0;
    output this_5_2_0_we0;
    output [63:0] this_5_2_0_d0;
    input [63:0] this_5_2_0_q0;
    output [2:0] this_5_2_1_address0;
    output this_5_2_1_ce0;
    output this_5_2_1_we0;
    output [63:0] this_5_2_1_d0;
    input [63:0] this_5_2_1_q0;
    output [2:0] this_5_2_2_address0;
    output this_5_2_2_ce0;
    output this_5_2_2_we0;
    output [63:0] this_5_2_2_d0;
    input [63:0] this_5_2_2_q0;
    output [2:0] this_5_2_3_address0;
    output this_5_2_3_ce0;
    output this_5_2_3_we0;
    output [63:0] this_5_2_3_d0;
    input [63:0] this_5_2_3_q0;
    output [2:0] this_5_3_0_address0;
    output this_5_3_0_ce0;
    output this_5_3_0_we0;
    output [63:0] this_5_3_0_d0;
    input [63:0] this_5_3_0_q0;
    output [2:0] this_5_3_1_address0;
    output this_5_3_1_ce0;
    output this_5_3_1_we0;
    output [63:0] this_5_3_1_d0;
    input [63:0] this_5_3_1_q0;
    output [2:0] this_5_3_2_address0;
    output this_5_3_2_ce0;
    output this_5_3_2_we0;
    output [63:0] this_5_3_2_d0;
    input [63:0] this_5_3_2_q0;
    output [2:0] this_5_3_3_address0;
    output this_5_3_3_ce0;
    output this_5_3_3_we0;
    output [63:0] this_5_3_3_d0;
    input [63:0] this_5_3_3_q0;
    output [2:0] this_6_0_0_address0;
    output this_6_0_0_ce0;
    output this_6_0_0_we0;
    output [63:0] this_6_0_0_d0;
    input [63:0] this_6_0_0_q0;
    output [2:0] this_6_0_1_address0;
    output this_6_0_1_ce0;
    output this_6_0_1_we0;
    output [63:0] this_6_0_1_d0;
    input [63:0] this_6_0_1_q0;
    output [2:0] this_6_0_2_address0;
    output this_6_0_2_ce0;
    output this_6_0_2_we0;
    output [63:0] this_6_0_2_d0;
    input [63:0] this_6_0_2_q0;
    output [2:0] this_6_0_3_address0;
    output this_6_0_3_ce0;
    output this_6_0_3_we0;
    output [63:0] this_6_0_3_d0;
    input [63:0] this_6_0_3_q0;
    output [2:0] this_6_1_0_address0;
    output this_6_1_0_ce0;
    output this_6_1_0_we0;
    output [63:0] this_6_1_0_d0;
    input [63:0] this_6_1_0_q0;
    output [2:0] this_6_1_1_address0;
    output this_6_1_1_ce0;
    output this_6_1_1_we0;
    output [63:0] this_6_1_1_d0;
    input [63:0] this_6_1_1_q0;
    output [2:0] this_6_1_2_address0;
    output this_6_1_2_ce0;
    output this_6_1_2_we0;
    output [63:0] this_6_1_2_d0;
    input [63:0] this_6_1_2_q0;
    output [2:0] this_6_1_3_address0;
    output this_6_1_3_ce0;
    output this_6_1_3_we0;
    output [63:0] this_6_1_3_d0;
    input [63:0] this_6_1_3_q0;
    output [2:0] this_6_2_0_address0;
    output this_6_2_0_ce0;
    output this_6_2_0_we0;
    output [63:0] this_6_2_0_d0;
    input [63:0] this_6_2_0_q0;
    output [2:0] this_6_2_1_address0;
    output this_6_2_1_ce0;
    output this_6_2_1_we0;
    output [63:0] this_6_2_1_d0;
    input [63:0] this_6_2_1_q0;
    output [2:0] this_6_2_2_address0;
    output this_6_2_2_ce0;
    output this_6_2_2_we0;
    output [63:0] this_6_2_2_d0;
    input [63:0] this_6_2_2_q0;
    output [2:0] this_6_2_3_address0;
    output this_6_2_3_ce0;
    output this_6_2_3_we0;
    output [63:0] this_6_2_3_d0;
    input [63:0] this_6_2_3_q0;
    output [2:0] this_6_3_0_address0;
    output this_6_3_0_ce0;
    output this_6_3_0_we0;
    output [63:0] this_6_3_0_d0;
    input [63:0] this_6_3_0_q0;
    output [2:0] this_6_3_1_address0;
    output this_6_3_1_ce0;
    output this_6_3_1_we0;
    output [63:0] this_6_3_1_d0;
    input [63:0] this_6_3_1_q0;
    output [2:0] this_6_3_2_address0;
    output this_6_3_2_ce0;
    output this_6_3_2_we0;
    output [63:0] this_6_3_2_d0;
    input [63:0] this_6_3_2_q0;
    output [2:0] this_6_3_3_address0;
    output this_6_3_3_ce0;
    output this_6_3_3_we0;
    output [63:0] this_6_3_3_d0;
    input [63:0] this_6_3_3_q0;
    output [2:0] this_7_address0;
    output this_7_ce0;
    output this_7_we0;
    output [63:0] this_7_d0;
    input [63:0] this_7_q0;
    input [63:0] p_read;
    input [63:0] p_read1;
    input [63:0] p_read2;
    input [63:0] p_read3;
    input [63:0] p_read4;
    input [63:0] p_read5;
    input [63:0] p_read6;
    input [63:0] p_read7;
    input [63:0] p_read8;
    input [63:0] p_read9;
    input [63:0] p_read10;
    input [63:0] p_read11;
    input [63:0] p_read12;
    input [63:0] p_read13;
    input [63:0] p_read14;
    input [63:0] p_read15;
    input [63:0] p_read16;
    input [63:0] p_read17;
    input [63:0] p_read18;
    input [63:0] p_read19;
    input [63:0] p_read20;
    input [63:0] p_read21;
    input [63:0] p_read22;
    input [63:0] p_read23;
    input [63:0] p_read24;
    input [63:0] p_read25;
    input [63:0] p_read26;
    input [63:0] p_read27;
    input [63:0] p_read28;
    input [63:0] p_read29;
    input [63:0] p_read30;
    input [63:0] p_read31;
    input [63:0] p_read32;
    input [63:0] p_read33;
    input [63:0] p_read34;
    input [63:0] p_read35;
    input [63:0] p_read36;
    input [63:0] p_read37;
    input [63:0] p_read38;
    input [63:0] p_read39;
    input [63:0] p_read40;
    input [63:0] p_read41;
    input [63:0] p_read42;
    input [63:0] p_read43;
    input [63:0] p_read44;
    input [63:0] p_read45;
    input [63:0] p_read46;
    input [63:0] p_read47;
    input [63:0] p_read48;
    input [63:0] p_read49;
    input [63:0] p_read50;
    input [63:0] p_read51;
    input [63:0] p_read52;
    input [63:0] p_read53;
    input [63:0] p_read54;
    input [63:0] p_read55;
    input [63:0] p_read56;
    input [63:0] p_read57;
    input [63:0] p_read58;
    input [63:0] p_read59;
    input [63:0] p_read60;
    input [63:0] p_read61;
    input [63:0] p_read62;
    input [63:0] p_read63;
    output [6:0] this_15_address0;
    output this_15_ce0;
    output this_15_we0;
    output [63:0] this_15_d0;
    input [63:0] this_15_q0;
    output [6:0] this_15_address1;
    output this_15_ce1;
    output this_15_we1;
    output [63:0] this_15_d1;
    input [63:0] this_15_q1;
    output [5:0] this_16_address0;
    output this_16_ce0;
    output this_16_we0;
    output [63:0] this_16_d0;
    input [63:0] this_16_q0;
    output [5:0] this_16_address1;
    output this_16_ce1;
    input [63:0] this_16_q1;
    input [63:0] l_TColl_0_0_0_constprop_i;
    output [63:0] l_TColl_0_0_0_constprop_o;
    output l_TColl_0_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_1_constprop_i;
    output [63:0] l_TColl_0_0_1_constprop_o;
    output l_TColl_0_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_2_constprop_i;
    output [63:0] l_TColl_0_0_2_constprop_o;
    output l_TColl_0_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_0_3_constprop_i;
    output [63:0] l_TColl_0_0_3_constprop_o;
    output l_TColl_0_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_0_constprop_i;
    output [63:0] l_TColl_1_0_0_constprop_o;
    output l_TColl_1_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_1_constprop_i;
    output [63:0] l_TColl_1_0_1_constprop_o;
    output l_TColl_1_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_2_constprop_i;
    output [63:0] l_TColl_1_0_2_constprop_o;
    output l_TColl_1_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_0_3_constprop_i;
    output [63:0] l_TColl_1_0_3_constprop_o;
    output l_TColl_1_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_0_constprop_i;
    output [63:0] l_TColl_2_0_0_constprop_o;
    output l_TColl_2_0_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_1_constprop_i;
    output [63:0] l_TColl_2_0_1_constprop_o;
    output l_TColl_2_0_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_2_constprop_i;
    output [63:0] l_TColl_2_0_2_constprop_o;
    output l_TColl_2_0_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_0_3_constprop_i;
    output [63:0] l_TColl_2_0_3_constprop_o;
    output l_TColl_2_0_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_0_constprop_i;
    output [63:0] l_TColl_0_1_0_constprop_o;
    output l_TColl_0_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_1_constprop_i;
    output [63:0] l_TColl_0_1_1_constprop_o;
    output l_TColl_0_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_2_constprop_i;
    output [63:0] l_TColl_0_1_2_constprop_o;
    output l_TColl_0_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_1_3_constprop_i;
    output [63:0] l_TColl_0_1_3_constprop_o;
    output l_TColl_0_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_0_constprop_i;
    output [63:0] l_TColl_1_1_0_constprop_o;
    output l_TColl_1_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_1_constprop_i;
    output [63:0] l_TColl_1_1_1_constprop_o;
    output l_TColl_1_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_2_constprop_i;
    output [63:0] l_TColl_1_1_2_constprop_o;
    output l_TColl_1_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_1_3_constprop_i;
    output [63:0] l_TColl_1_1_3_constprop_o;
    output l_TColl_1_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_0_constprop_i;
    output [63:0] l_TColl_2_1_0_constprop_o;
    output l_TColl_2_1_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_1_constprop_i;
    output [63:0] l_TColl_2_1_1_constprop_o;
    output l_TColl_2_1_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_2_constprop_i;
    output [63:0] l_TColl_2_1_2_constprop_o;
    output l_TColl_2_1_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_1_3_constprop_i;
    output [63:0] l_TColl_2_1_3_constprop_o;
    output l_TColl_2_1_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_0_constprop_i;
    output [63:0] l_TColl_0_2_0_constprop_o;
    output l_TColl_0_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_1_constprop_i;
    output [63:0] l_TColl_0_2_1_constprop_o;
    output l_TColl_0_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_2_constprop_i;
    output [63:0] l_TColl_0_2_2_constprop_o;
    output l_TColl_0_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_2_3_constprop_i;
    output [63:0] l_TColl_0_2_3_constprop_o;
    output l_TColl_0_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_0_constprop_i;
    output [63:0] l_TColl_1_2_0_constprop_o;
    output l_TColl_1_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_1_constprop_i;
    output [63:0] l_TColl_1_2_1_constprop_o;
    output l_TColl_1_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_2_constprop_i;
    output [63:0] l_TColl_1_2_2_constprop_o;
    output l_TColl_1_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_2_3_constprop_i;
    output [63:0] l_TColl_1_2_3_constprop_o;
    output l_TColl_1_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_0_constprop_i;
    output [63:0] l_TColl_2_2_0_constprop_o;
    output l_TColl_2_2_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_1_constprop_i;
    output [63:0] l_TColl_2_2_1_constprop_o;
    output l_TColl_2_2_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_2_constprop_i;
    output [63:0] l_TColl_2_2_2_constprop_o;
    output l_TColl_2_2_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_2_3_constprop_i;
    output [63:0] l_TColl_2_2_3_constprop_o;
    output l_TColl_2_2_3_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_0_constprop_i;
    output [63:0] l_TColl_0_3_0_constprop_o;
    output l_TColl_0_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_1_constprop_i;
    output [63:0] l_TColl_0_3_1_constprop_o;
    output l_TColl_0_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_2_constprop_i;
    output [63:0] l_TColl_0_3_2_constprop_o;
    output l_TColl_0_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_0_3_3_constprop_i;
    output [63:0] l_TColl_0_3_3_constprop_o;
    output l_TColl_0_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_0_constprop_i;
    output [63:0] l_TColl_1_3_0_constprop_o;
    output l_TColl_1_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_1_constprop_i;
    output [63:0] l_TColl_1_3_1_constprop_o;
    output l_TColl_1_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_2_constprop_i;
    output [63:0] l_TColl_1_3_2_constprop_o;
    output l_TColl_1_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_1_3_3_constprop_i;
    output [63:0] l_TColl_1_3_3_constprop_o;
    output l_TColl_1_3_3_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_0_constprop_i;
    output [63:0] l_TColl_2_3_0_constprop_o;
    output l_TColl_2_3_0_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_1_constprop_i;
    output [63:0] l_TColl_2_3_1_constprop_o;
    output l_TColl_2_3_1_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_2_constprop_i;
    output [63:0] l_TColl_2_3_2_constprop_o;
    output l_TColl_2_3_2_constprop_o_ap_vld;
    input [63:0] l_TColl_2_3_3_constprop_i;
    output [63:0] l_TColl_2_3_3_constprop_o;
    output l_TColl_2_3_3_constprop_o_ap_vld;
    output [63:0] grp_fu_2427_p_din0;
    output [63:0] grp_fu_2427_p_din1;
    output [0:0] grp_fu_2427_p_opcode;
    input [63:0] grp_fu_2427_p_dout0;
    output grp_fu_2427_p_ce;
    output [63:0] grp_fu_2403_p_din0;
    output [63:0] grp_fu_2403_p_din1;
    output [1:0] grp_fu_2403_p_opcode;
    input [63:0] grp_fu_2403_p_dout0;
    output grp_fu_2403_p_ce;
    output [63:0] grp_fu_2431_p_din0;
    output [63:0] grp_fu_2431_p_din1;
    input [63:0] grp_fu_2431_p_dout0;
    output grp_fu_2431_p_ce;
    output [63:0] grp_fu_2407_p_din0;
    output [63:0] grp_fu_2407_p_din1;
    output [1:0] grp_fu_2407_p_opcode;
    input [63:0] grp_fu_2407_p_dout0;
    output grp_fu_2407_p_ce;
    output [63:0] grp_fu_2411_p_din0;
    output [63:0] grp_fu_2411_p_din1;
    output [1:0] grp_fu_2411_p_opcode;
    input [63:0] grp_fu_2411_p_dout0;
    output grp_fu_2411_p_ce;
    output [63:0] grp_fu_2415_p_din0;
    output [63:0] grp_fu_2415_p_din1;
    output [1:0] grp_fu_2415_p_opcode;
    input [63:0] grp_fu_2415_p_dout0;
    output grp_fu_2415_p_ce;
    output [63:0] grp_fu_2419_p_din0;
    output [63:0] grp_fu_2419_p_din1;
    output [1:0] grp_fu_2419_p_opcode;
    input [63:0] grp_fu_2419_p_dout0;
    output grp_fu_2419_p_ce;
    output [63:0] grp_fu_2423_p_din0;
    output [63:0] grp_fu_2423_p_din1;
    output [1:0] grp_fu_2423_p_opcode;
    input [63:0] grp_fu_2423_p_dout0;
    output grp_fu_2423_p_ce;
    output [63:0] grp_fu_2435_p_din0;
    output [63:0] grp_fu_2435_p_din1;
    input [63:0] grp_fu_2435_p_dout0;
    output grp_fu_2435_p_ce;
    output [63:0] grp_fu_2439_p_din0;
    output [63:0] grp_fu_2439_p_din1;
    input [63:0] grp_fu_2439_p_dout0;
    output grp_fu_2439_p_ce;
    output [63:0] grp_fu_2443_p_din0;
    output [63:0] grp_fu_2443_p_din1;
    input [63:0] grp_fu_2443_p_dout0;
    output grp_fu_2443_p_ce;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg [63:0] l_TColl_0_0_0_constprop_o;
    reg [63:0] l_TColl_0_0_1_constprop_o;
    reg [63:0] l_TColl_0_0_2_constprop_o;
    reg [63:0] l_TColl_0_0_3_constprop_o;
    reg [63:0] l_TColl_1_0_0_constprop_o;
    reg [63:0] l_TColl_1_0_1_constprop_o;
    reg [63:0] l_TColl_1_0_2_constprop_o;
    reg [63:0] l_TColl_1_0_3_constprop_o;
    reg [63:0] l_TColl_2_0_0_constprop_o;
    reg [63:0] l_TColl_2_0_1_constprop_o;
    reg [63:0] l_TColl_2_0_2_constprop_o;
    reg [63:0] l_TColl_2_0_3_constprop_o;
    reg [63:0] l_TColl_0_1_0_constprop_o;
    reg [63:0] l_TColl_0_1_1_constprop_o;
    reg [63:0] l_TColl_0_1_2_constprop_o;
    reg [63:0] l_TColl_0_1_3_constprop_o;
    reg [63:0] l_TColl_1_1_0_constprop_o;
    reg [63:0] l_TColl_1_1_1_constprop_o;
    reg [63:0] l_TColl_1_1_2_constprop_o;
    reg [63:0] l_TColl_1_1_3_constprop_o;
    reg [63:0] l_TColl_2_1_0_constprop_o;
    reg [63:0] l_TColl_2_1_1_constprop_o;
    reg [63:0] l_TColl_2_1_2_constprop_o;
    reg [63:0] l_TColl_2_1_3_constprop_o;
    reg [63:0] l_TColl_0_2_0_constprop_o;
    reg [63:0] l_TColl_0_2_1_constprop_o;
    reg [63:0] l_TColl_0_2_2_constprop_o;
    reg [63:0] l_TColl_0_2_3_constprop_o;
    reg [63:0] l_TColl_1_2_0_constprop_o;
    reg [63:0] l_TColl_1_2_1_constprop_o;
    reg [63:0] l_TColl_1_2_2_constprop_o;
    reg [63:0] l_TColl_1_2_3_constprop_o;
    reg [63:0] l_TColl_2_2_0_constprop_o;
    reg [63:0] l_TColl_2_2_1_constprop_o;
    reg [63:0] l_TColl_2_2_2_constprop_o;
    reg [63:0] l_TColl_2_2_3_constprop_o;
    reg [63:0] l_TColl_0_3_0_constprop_o;
    reg [63:0] l_TColl_0_3_1_constprop_o;
    reg [63:0] l_TColl_0_3_2_constprop_o;
    reg [63:0] l_TColl_0_3_3_constprop_o;
    reg [63:0] l_TColl_1_3_0_constprop_o;
    reg [63:0] l_TColl_1_3_1_constprop_o;
    reg [63:0] l_TColl_1_3_2_constprop_o;
    reg [63:0] l_TColl_1_3_3_constprop_o;
    reg [63:0] l_TColl_2_3_0_constprop_o;
    reg [63:0] l_TColl_2_3_1_constprop_o;
    reg [63:0] l_TColl_2_3_2_constprop_o;
    reg [63:0] l_TColl_2_3_3_constprop_o;

    (* fsm_encoding = "none" *) reg [337:0] ap_CS_fsm;
    wire ap_CS_fsm_state1;
    reg [15:0] lfsr;
    reg [2:0] goal_address0;
    reg goal_ce0;
    wire [63:0] goal_q0;
    wire [63:0] grp_fu_1462_p2;
    reg [63:0] reg_1470;
    wire ap_CS_fsm_state79;
    wire ap_CS_fsm_state142;
    wire ap_CS_fsm_state274;
    wire ap_CS_fsm_state335;
    wire ap_CS_fsm_state2;
    reg [31:0] numVertices_1_reg_2362;
    wire ap_CS_fsm_state3;
    wire [11:0] trunc_ln83_fu_1483_p1;
    reg [11:0] trunc_ln83_reg_2369;
    wire [9:0] trunc_ln83_1_fu_1487_p1;
    reg [9:0] trunc_ln83_1_reg_2374;
    wire [0:0] icmp_ln107_fu_1491_p2;
    reg [0:0] icmp_ln107_reg_2379;
    reg [14:0] lshr_ln_reg_2386;
    wire ap_CS_fsm_state5;
    wire [0:0] xor_ln38_fu_1558_p2;
    reg [0:0] xor_ln38_reg_2391;
    wire [31:0] zext_ln47_fu_1576_p1;
    wire ap_CS_fsm_state6;
    wire [31:0] grp_fu_1436_p1;
    reg [31:0] conv_i1_reg_2401;
    wire ap_CS_fsm_state11;
    wire [31:0] grp_fu_1431_p2;
    reg [31:0] div_i_reg_2406;
    wire ap_CS_fsm_state15;
    wire [63:0] grp_fu_1439_p1;
    reg [63:0] conv_reg_2411;
    wire ap_CS_fsm_state17;
    wire [0:0] icmp_ln110_fu_1598_p2;
    reg [0:0] icmp_ln110_reg_2417;
    wire ap_CS_fsm_state18;
    wire [0:0] icmp_ln110_1_fu_1604_p2;
    reg [0:0] icmp_ln110_1_reg_2422;
    wire [0:0] and_ln110_fu_1614_p2;
    reg [0:0] and_ln110_reg_2427;
    wire ap_CS_fsm_state19;
    wire [12:0] sub_ln130_fu_1634_p2;
    reg [12:0] sub_ln130_reg_2431;
    wire ap_CS_fsm_state20;
    wire [31:0] select_ln96_fu_1664_p3;
    reg [31:0] select_ln96_reg_2439;
    wire [34:0] sub_ln296_fu_1690_p2;
    reg [34:0] sub_ln296_reg_2445;
    wire ap_CS_fsm_state80;
    wire [12:0] sub_ln114_fu_1720_p2;
    reg [12:0] sub_ln114_reg_2450;
    wire ap_CS_fsm_state82;
    wire [0:0] and_ln119_fu_1767_p2;
    reg [0:0] and_ln119_reg_2458;
    wire ap_CS_fsm_state144;
    wire [63:0] grp_fu_1448_p2;
    reg [63:0] f_reg_2462;
    wire ap_CS_fsm_state203;
    wire [0:0] and_ln188_fu_1809_p2;
    reg [0:0] and_ln188_reg_2467;
    wire ap_CS_fsm_state206;
    wire ap_CS_fsm_state215;
    wire [11:0] trunc_ln83_2_fu_1829_p1;
    reg [11:0] trunc_ln83_2_reg_2482;
    wire [9:0] trunc_ln83_3_fu_1833_p1;
    reg [9:0] trunc_ln83_3_reg_2487;
    wire [31:0] select_ln96_5_fu_1859_p3;
    reg [31:0] select_ln96_5_reg_2492;
    wire [34:0] sub_ln296_1_fu_1885_p2;
    reg [34:0] sub_ln296_1_reg_2498;
    wire ap_CS_fsm_state275;
    wire [12:0] sub_ln294_fu_1915_p2;
    reg [12:0] sub_ln294_reg_2503;
    wire ap_CS_fsm_state277;
    wire [0:0] icmp_ln138_fu_1944_p2;
    reg [0:0] icmp_ln138_reg_2511;
    wire ap_CS_fsm_state336;
    wire [0:0] icmp_ln138_1_fu_1950_p2;
    reg [0:0] icmp_ln138_1_reg_2516;
    wire [12:0] sub_ln139_fu_1980_p2;
    reg [12:0] sub_ln139_reg_2524;
    wire ap_CS_fsm_state337;
    reg [2:0] ang_address0;
    reg ang_ce0;
    reg ang_we0;
    wire [63:0] ang_q0;
    reg [12:0] rrtVertices_address0;
    reg rrtVertices_ce0;
    reg rrtVertices_we0;
    reg [63:0] rrtVertices_d0;
    wire [63:0] rrtVertices_q0;
    reg [2:0] qRand_address0;
    reg qRand_ce0;
    reg qRand_we0;
    reg [63:0] qRand_d0;
    wire [63:0] qRand_q0;
    reg [2:0] qNear_address0;
    reg qNear_ce0;
    reg qNear_we0;
    wire [63:0] qNear_q0;
    reg [2:0] qConnect_address0;
    reg qConnect_ce0;
    reg qConnect_we0;
    reg [63:0] qConnect_d0;
    wire [63:0] qConnect_q0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_d0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_d0;
    wire [15:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out_ap_vld;
    wire [5:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out_ap_vld;
    wire [31:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din0;
    wire [31:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_ce;
    wire [31:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_din0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_ce;
    wire [31:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_din0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din1;
    wire [0:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_d0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_dist_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_dist_out_ap_vld;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_ce0;
    wire [11:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out_ap_vld;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din1;
    wire [4:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_d0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_dist_4_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_dist_4_out_ap_vld;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_d0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_d0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din1;
    wire [0:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din1;
    wire [0:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_ready;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_ce0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_d0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din1;
    wire [0:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din1;
    wire [0:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_d0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_ce0;
    wire grp_detectCollNode_fu_1055_ap_start;
    wire grp_detectCollNode_fu_1055_ap_done;
    wire grp_detectCollNode_fu_1055_ap_idle;
    wire grp_detectCollNode_fu_1055_ap_ready;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_0_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_0_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_0_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_0_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_0_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_0_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_1_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_1_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_1_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_1_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_1_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_1_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_2_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_2_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_2_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_2_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_2_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_2_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_3_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_3_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_3_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_3_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_3_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_3_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_4_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_4_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_4_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_4_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_4_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_4_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_5_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_5_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_5_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_5_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_5_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_5_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_6_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_6_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_6_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_6_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_6_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_6_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_7_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_7_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_7_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_7_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_7_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_7_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_8_0_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_8_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_8_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_8_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_env_0_8_2_address0;
    wire grp_detectCollNode_fu_1055_this_env_0_8_2_ce0;
    wire [6:0] grp_detectCollNode_fu_1055_this_env_1_address0;
    wire grp_detectCollNode_fu_1055_this_env_1_ce0;
    wire [6:0] grp_detectCollNode_fu_1055_this_env_1_address1;
    wire grp_detectCollNode_fu_1055_this_env_1_ce1;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_0_0_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_0_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_0_1_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_0_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_0_2_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_0_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_0_3_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_0_3_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_1_0_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_1_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_1_1_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_1_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_1_2_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_1_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_1_3_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_1_3_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_2_0_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_2_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_2_1_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_2_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_2_2_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_2_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_2_3_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_2_3_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_3_0_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_3_0_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_3_1_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_3_1_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_3_2_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_3_2_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TLink_3_3_address0;
    wire grp_detectCollNode_fu_1055_this_TLink_3_3_ce0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_0_0_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_0_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_0_1_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_0_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_0_2_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_0_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_0_3_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_0_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_0_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_1_0_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_1_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_1_1_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_1_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_1_2_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_1_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_1_3_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_1_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_1_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_2_0_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_2_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_2_1_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_2_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_2_2_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_2_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_2_3_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_2_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_2_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_3_0_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_3_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_3_1_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_3_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_3_2_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_3_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TJoint_3_3_address0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TJoint_3_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TJoint_3_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_0_0_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_0_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_0_1_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_0_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_0_2_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_0_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_0_3_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_0_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_0_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_1_0_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_1_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_1_1_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_1_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_1_2_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_1_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_1_3_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_1_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_1_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_2_0_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_2_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_2_1_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_2_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_2_2_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_2_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_2_3_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_2_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_2_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_3_0_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_0_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_0_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_3_0_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_3_1_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_1_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_1_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_3_1_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_3_2_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_2_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_2_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_3_2_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_TCurr_3_3_address0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_3_ce0;
    wire grp_detectCollNode_fu_1055_this_TCurr_3_3_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_TCurr_3_3_d0;
    wire [2:0] grp_detectCollNode_fu_1055_this_q_address0;
    wire grp_detectCollNode_fu_1055_this_q_ce0;
    wire grp_detectCollNode_fu_1055_this_q_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_q_d0;
    wire [6:0] grp_detectCollNode_fu_1055_this_cPoints_address0;
    wire grp_detectCollNode_fu_1055_this_cPoints_ce0;
    wire grp_detectCollNode_fu_1055_this_cPoints_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_cPoints_d0;
    wire [6:0] grp_detectCollNode_fu_1055_this_cPoints_address1;
    wire grp_detectCollNode_fu_1055_this_cPoints_ce1;
    wire grp_detectCollNode_fu_1055_this_cPoints_we1;
    wire [63:0] grp_detectCollNode_fu_1055_this_cPoints_d1;
    wire [5:0] grp_detectCollNode_fu_1055_this_cAxes_address0;
    wire grp_detectCollNode_fu_1055_this_cAxes_ce0;
    wire grp_detectCollNode_fu_1055_this_cAxes_we0;
    wire [63:0] grp_detectCollNode_fu_1055_this_cAxes_d0;
    wire [5:0] grp_detectCollNode_fu_1055_this_cAxes_address1;
    wire grp_detectCollNode_fu_1055_this_cAxes_ce1;
    wire [2:0] grp_detectCollNode_fu_1055_ang_address0;
    wire grp_detectCollNode_fu_1055_ang_ce0;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o_ap_vld;
    wire [63:0] grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o;
    wire grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o_ap_vld;
    wire [0:0] grp_detectCollNode_fu_1055_ap_return;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2529_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2529_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2529_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2529_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2533_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2533_p_din1;
    wire grp_detectCollNode_fu_1055_grp_fu_2533_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2537_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2537_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2537_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2537_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2541_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2541_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2541_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2541_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2545_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2545_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2545_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2545_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2549_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2549_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2549_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2549_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2553_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2553_p_din1;
    wire [1:0] grp_detectCollNode_fu_1055_grp_fu_2553_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_2553_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2557_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2557_p_din1;
    wire grp_detectCollNode_fu_1055_grp_fu_2557_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2561_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2561_p_din1;
    wire grp_detectCollNode_fu_1055_grp_fu_2561_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2565_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_2565_p_din1;
    wire grp_detectCollNode_fu_1055_grp_fu_2565_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_1454_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_1454_p_din1;
    wire [4:0] grp_detectCollNode_fu_1055_grp_fu_1454_p_opcode;
    wire grp_detectCollNode_fu_1055_grp_fu_1454_p_ce;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_1462_p_din0;
    wire [63:0] grp_detectCollNode_fu_1055_grp_fu_1462_p_din1;
    wire grp_detectCollNode_fu_1055_grp_fu_1462_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_dist_6_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_dist_6_out_ap_vld;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_ready;
    wire   [12:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_ce0;
    wire [11:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out_ap_vld;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din1;
    wire [4:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_dist_10_out;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_dist_10_out_ap_vld;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_ce0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din1;
    wire [1:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_opcode;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_ce;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din1;
    wire grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_ce;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_done;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_idle;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_ready;
    wire [12:0] grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_ce0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_we0;
    wire [63:0] grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_d0;
    wire [2:0] grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_address0;
    wire grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_ce0;
    reg [63:0] s_reg_960;
    wire ap_CS_fsm_state204;
    reg ap_block_state204_on_subcall_done;
    reg grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg;
    reg grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg;
    wire ap_CS_fsm_state4;
    reg grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg;
    reg grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg;
    wire ap_CS_fsm_state21;
    wire ap_CS_fsm_state22;
    reg grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg;
    wire ap_CS_fsm_state81;
    reg [11:0] bestIdx_3_loc_fu_540;
    reg grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg;
    wire ap_CS_fsm_state83;
    reg grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg;
    wire ap_CS_fsm_state84;
    wire ap_CS_fsm_state85;
    reg grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg;
    wire ap_CS_fsm_state145;
    reg grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg;
    reg grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg;
    wire ap_CS_fsm_state207;
    reg grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg;
    wire ap_CS_fsm_state216;
    reg grp_detectCollNode_fu_1055_ap_start_reg;
    wire ap_CS_fsm_state208;
    wire ap_CS_fsm_state209;
    reg grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg;
    reg ap_block_state209_on_subcall_done;
    wire ap_CS_fsm_state217;
    reg grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg;
    wire ap_CS_fsm_state276;
    reg [11:0] bestIdx_6_loc_fu_528;
    reg grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg;
    wire ap_CS_fsm_state278;
    reg grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg;
    wire [0:0] and_ln138_fu_1960_p2;
    wire ap_CS_fsm_state338;
    wire [15:0] rand_int_fu_1564_p3;
    reg [31:0] numVertices_fu_520;
    wire [31:0] numVertices_2_fu_1815_p2;
    wire ap_CS_fsm_state279;
    wire ap_CS_fsm_state218;
    wire ap_CS_fsm_state86;
    wire ap_CS_fsm_state23;
    reg [31:0] grp_fu_1431_p0;
    reg [31:0] grp_fu_1431_p1;
    wire ap_CS_fsm_state12;
    reg [31:0] grp_fu_1436_p0;
    reg [31:0] grp_fu_1439_p0;
    wire ap_CS_fsm_state16;
    reg [63:0] grp_fu_1454_p0;
    reg [63:0] grp_fu_1454_p1;
    wire ap_CS_fsm_state143;
    wire ap_CS_fsm_state205;
    reg [63:0] grp_fu_1462_p1;
    wire [0:0] tmp_16_fu_1512_p3;
    wire [0:0] trunc_ln37_fu_1508_p1;
    wire [0:0] tmp_17_fu_1520_p3;
    wire [0:0] tmp_18_fu_1528_p3;
    wire [0:0] xor_ln38_3_fu_1552_p2;
    wire [0:0] xor_ln38_2_fu_1546_p2;
    wire [63:0] bitcast_ln110_fu_1581_p1;
    wire [10:0] tmp_262_fu_1584_p4;
    wire [51:0] trunc_ln110_fu_1594_p1;
    wire [0:0] or_ln110_fu_1610_p2;
    wire [0:0] grp_fu_1454_p2;
    wire [12:0] tmp_fu_1620_p3;
    wire [12:0] tmp_24_fu_1627_p3;
    wire [30:0] tmp_19_fu_1644_p4;
    wire [0:0] icmp_fu_1653_p2;
    wire [31:0] add_ln96_2_fu_1659_p2;
    wire [32:0] tmp_25_fu_1679_p3;
    wire [34:0] p_shl_fu_1672_p3;
    wire [34:0] zext_ln296_fu_1686_p1;
    wire [9:0] empty_fu_1700_p1;
    wire [12:0] tmp_26_fu_1704_p3;
    wire [12:0] tmp_27_fu_1712_p3;
    wire [63:0] bitcast_ln119_fu_1731_p1;
    wire [10:0] tmp_264_fu_1735_p4;
    wire [51:0] trunc_ln119_fu_1745_p1;
    wire [0:0] icmp_ln119_1_fu_1755_p2;
    wire [0:0] icmp_ln119_fu_1749_p2;
    wire [0:0] or_ln119_fu_1761_p2;
    wire [63:0] bitcast_ln188_fu_1773_p1;
    wire [10:0] tmp_266_fu_1777_p4;
    wire [51:0] trunc_ln188_fu_1787_p1;
    wire [0:0] icmp_ln188_1_fu_1797_p2;
    wire [0:0] icmp_ln188_fu_1791_p2;
    wire [0:0] or_ln188_fu_1803_p2;
    wire [30:0] tmp_20_fu_1837_p4;
    wire [0:0] icmp35_fu_1847_p2;
    wire [31:0] add_ln96_fu_1853_p2;
    wire [32:0] tmp_30_fu_1874_p3;
    wire [34:0] p_shl1_fu_1867_p3;
    wire [34:0] zext_ln296_1_fu_1881_p1;
    wire [9:0] empty_64_fu_1895_p1;
    wire [12:0] tmp_31_fu_1899_p3;
    wire [12:0] tmp_32_fu_1907_p3;
    wire [63:0] bitcast_ln138_fu_1926_p1;
    wire [10:0] tmp_268_fu_1930_p4;
    wire [51:0] trunc_ln138_fu_1940_p1;
    wire [0:0] or_ln138_fu_1956_p2;
    wire [12:0] tmp_35_fu_1966_p3;
    wire [12:0] tmp_36_fu_1973_p3;
    reg grp_fu_1431_ce;
    reg grp_fu_1436_ce;
    reg grp_fu_1439_ce;
    reg grp_fu_1442_ce;
    wire ap_CS_fsm_state210;
    wire ap_CS_fsm_state211;
    wire ap_CS_fsm_state212;
    wire ap_CS_fsm_state213;
    wire ap_CS_fsm_state214;
    reg grp_fu_1454_ce;
    reg [4:0] grp_fu_1454_opcode;
    reg [63:0] grp_fu_1462_p0;
    reg grp_fu_1462_ce;
    reg [63:0] grp_fu_2529_p0;
    reg [63:0] grp_fu_2529_p1;
    reg [1:0] grp_fu_2529_opcode;
    reg grp_fu_2529_ce;
    reg [63:0] grp_fu_2533_p0;
    reg [63:0] grp_fu_2533_p1;
    reg grp_fu_2533_ce;
    reg [63:0] grp_fu_2537_p0;
    reg [63:0] grp_fu_2537_p1;
    reg [1:0] grp_fu_2537_opcode;
    reg grp_fu_2537_ce;
    reg grp_fu_2541_ce;
    reg grp_fu_2545_ce;
    reg grp_fu_2549_ce;
    reg grp_fu_2553_ce;
    reg grp_fu_2557_ce;
    reg grp_fu_2561_ce;
    reg grp_fu_2565_ce;
    reg ap_block_state338_on_subcall_done;
    reg [337:0] ap_NS_fsm;
    reg ap_ST_fsm_state1_blk;
    reg ap_ST_fsm_state2_blk;
    wire ap_ST_fsm_state3_blk;
    reg ap_ST_fsm_state4_blk;
    wire ap_ST_fsm_state5_blk;
    wire ap_ST_fsm_state6_blk;
    wire ap_ST_fsm_state7_blk;
    wire ap_ST_fsm_state8_blk;
    wire ap_ST_fsm_state9_blk;
    wire ap_ST_fsm_state10_blk;
    wire ap_ST_fsm_state11_blk;
    wire ap_ST_fsm_state12_blk;
    wire ap_ST_fsm_state13_blk;
    wire ap_ST_fsm_state14_blk;
    wire ap_ST_fsm_state15_blk;
    wire ap_ST_fsm_state16_blk;
    wire ap_ST_fsm_state17_blk;
    wire ap_ST_fsm_state18_blk;
    wire ap_ST_fsm_state19_blk;
    reg ap_block_state20_on_subcall_done;
    reg ap_ST_fsm_state20_blk;
    wire ap_ST_fsm_state21_blk;
    reg ap_ST_fsm_state22_blk;
    wire ap_ST_fsm_state23_blk;
    wire ap_ST_fsm_state24_blk;
    wire ap_ST_fsm_state25_blk;
    wire ap_ST_fsm_state26_blk;
    wire ap_ST_fsm_state27_blk;
    wire ap_ST_fsm_state28_blk;
    wire ap_ST_fsm_state29_blk;
    wire ap_ST_fsm_state30_blk;
    wire ap_ST_fsm_state31_blk;
    wire ap_ST_fsm_state32_blk;
    wire ap_ST_fsm_state33_blk;
    wire ap_ST_fsm_state34_blk;
    wire ap_ST_fsm_state35_blk;
    wire ap_ST_fsm_state36_blk;
    wire ap_ST_fsm_state37_blk;
    wire ap_ST_fsm_state38_blk;
    wire ap_ST_fsm_state39_blk;
    wire ap_ST_fsm_state40_blk;
    wire ap_ST_fsm_state41_blk;
    wire ap_ST_fsm_state42_blk;
    wire ap_ST_fsm_state43_blk;
    wire ap_ST_fsm_state44_blk;
    wire ap_ST_fsm_state45_blk;
    wire ap_ST_fsm_state46_blk;
    wire ap_ST_fsm_state47_blk;
    wire ap_ST_fsm_state48_blk;
    wire ap_ST_fsm_state49_blk;
    wire ap_ST_fsm_state50_blk;
    wire ap_ST_fsm_state51_blk;
    wire ap_ST_fsm_state52_blk;
    wire ap_ST_fsm_state53_blk;
    wire ap_ST_fsm_state54_blk;
    wire ap_ST_fsm_state55_blk;
    wire ap_ST_fsm_state56_blk;
    wire ap_ST_fsm_state57_blk;
    wire ap_ST_fsm_state58_blk;
    wire ap_ST_fsm_state59_blk;
    wire ap_ST_fsm_state60_blk;
    wire ap_ST_fsm_state61_blk;
    wire ap_ST_fsm_state62_blk;
    wire ap_ST_fsm_state63_blk;
    wire ap_ST_fsm_state64_blk;
    wire ap_ST_fsm_state65_blk;
    wire ap_ST_fsm_state66_blk;
    wire ap_ST_fsm_state67_blk;
    wire ap_ST_fsm_state68_blk;
    wire ap_ST_fsm_state69_blk;
    wire ap_ST_fsm_state70_blk;
    wire ap_ST_fsm_state71_blk;
    wire ap_ST_fsm_state72_blk;
    wire ap_ST_fsm_state73_blk;
    wire ap_ST_fsm_state74_blk;
    wire ap_ST_fsm_state75_blk;
    wire ap_ST_fsm_state76_blk;
    wire ap_ST_fsm_state77_blk;
    wire ap_ST_fsm_state78_blk;
    wire ap_ST_fsm_state79_blk;
    wire ap_ST_fsm_state80_blk;
    reg ap_ST_fsm_state81_blk;
    wire ap_ST_fsm_state82_blk;
    reg ap_ST_fsm_state83_blk;
    wire ap_ST_fsm_state84_blk;
    reg ap_ST_fsm_state85_blk;
    wire ap_ST_fsm_state86_blk;
    wire ap_ST_fsm_state87_blk;
    wire ap_ST_fsm_state88_blk;
    wire ap_ST_fsm_state89_blk;
    wire ap_ST_fsm_state90_blk;
    wire ap_ST_fsm_state91_blk;
    wire ap_ST_fsm_state92_blk;
    wire ap_ST_fsm_state93_blk;
    wire ap_ST_fsm_state94_blk;
    wire ap_ST_fsm_state95_blk;
    wire ap_ST_fsm_state96_blk;
    wire ap_ST_fsm_state97_blk;
    wire ap_ST_fsm_state98_blk;
    wire ap_ST_fsm_state99_blk;
    wire ap_ST_fsm_state100_blk;
    wire ap_ST_fsm_state101_blk;
    wire ap_ST_fsm_state102_blk;
    wire ap_ST_fsm_state103_blk;
    wire ap_ST_fsm_state104_blk;
    wire ap_ST_fsm_state105_blk;
    wire ap_ST_fsm_state106_blk;
    wire ap_ST_fsm_state107_blk;
    wire ap_ST_fsm_state108_blk;
    wire ap_ST_fsm_state109_blk;
    wire ap_ST_fsm_state110_blk;
    wire ap_ST_fsm_state111_blk;
    wire ap_ST_fsm_state112_blk;
    wire ap_ST_fsm_state113_blk;
    wire ap_ST_fsm_state114_blk;
    wire ap_ST_fsm_state115_blk;
    wire ap_ST_fsm_state116_blk;
    wire ap_ST_fsm_state117_blk;
    wire ap_ST_fsm_state118_blk;
    wire ap_ST_fsm_state119_blk;
    wire ap_ST_fsm_state120_blk;
    wire ap_ST_fsm_state121_blk;
    wire ap_ST_fsm_state122_blk;
    wire ap_ST_fsm_state123_blk;
    wire ap_ST_fsm_state124_blk;
    wire ap_ST_fsm_state125_blk;
    wire ap_ST_fsm_state126_blk;
    wire ap_ST_fsm_state127_blk;
    wire ap_ST_fsm_state128_blk;
    wire ap_ST_fsm_state129_blk;
    wire ap_ST_fsm_state130_blk;
    wire ap_ST_fsm_state131_blk;
    wire ap_ST_fsm_state132_blk;
    wire ap_ST_fsm_state133_blk;
    wire ap_ST_fsm_state134_blk;
    wire ap_ST_fsm_state135_blk;
    wire ap_ST_fsm_state136_blk;
    wire ap_ST_fsm_state137_blk;
    wire ap_ST_fsm_state138_blk;
    wire ap_ST_fsm_state139_blk;
    wire ap_ST_fsm_state140_blk;
    wire ap_ST_fsm_state141_blk;
    wire ap_ST_fsm_state142_blk;
    wire ap_ST_fsm_state143_blk;
    wire ap_ST_fsm_state144_blk;
    reg ap_ST_fsm_state145_blk;
    wire ap_ST_fsm_state146_blk;
    wire ap_ST_fsm_state147_blk;
    wire ap_ST_fsm_state148_blk;
    wire ap_ST_fsm_state149_blk;
    wire ap_ST_fsm_state150_blk;
    wire ap_ST_fsm_state151_blk;
    wire ap_ST_fsm_state152_blk;
    wire ap_ST_fsm_state153_blk;
    wire ap_ST_fsm_state154_blk;
    wire ap_ST_fsm_state155_blk;
    wire ap_ST_fsm_state156_blk;
    wire ap_ST_fsm_state157_blk;
    wire ap_ST_fsm_state158_blk;
    wire ap_ST_fsm_state159_blk;
    wire ap_ST_fsm_state160_blk;
    wire ap_ST_fsm_state161_blk;
    wire ap_ST_fsm_state162_blk;
    wire ap_ST_fsm_state163_blk;
    wire ap_ST_fsm_state164_blk;
    wire ap_ST_fsm_state165_blk;
    wire ap_ST_fsm_state166_blk;
    wire ap_ST_fsm_state167_blk;
    wire ap_ST_fsm_state168_blk;
    wire ap_ST_fsm_state169_blk;
    wire ap_ST_fsm_state170_blk;
    wire ap_ST_fsm_state171_blk;
    wire ap_ST_fsm_state172_blk;
    wire ap_ST_fsm_state173_blk;
    wire ap_ST_fsm_state174_blk;
    wire ap_ST_fsm_state175_blk;
    wire ap_ST_fsm_state176_blk;
    wire ap_ST_fsm_state177_blk;
    wire ap_ST_fsm_state178_blk;
    wire ap_ST_fsm_state179_blk;
    wire ap_ST_fsm_state180_blk;
    wire ap_ST_fsm_state181_blk;
    wire ap_ST_fsm_state182_blk;
    wire ap_ST_fsm_state183_blk;
    wire ap_ST_fsm_state184_blk;
    wire ap_ST_fsm_state185_blk;
    wire ap_ST_fsm_state186_blk;
    wire ap_ST_fsm_state187_blk;
    wire ap_ST_fsm_state188_blk;
    wire ap_ST_fsm_state189_blk;
    wire ap_ST_fsm_state190_blk;
    wire ap_ST_fsm_state191_blk;
    wire ap_ST_fsm_state192_blk;
    wire ap_ST_fsm_state193_blk;
    wire ap_ST_fsm_state194_blk;
    wire ap_ST_fsm_state195_blk;
    wire ap_ST_fsm_state196_blk;
    wire ap_ST_fsm_state197_blk;
    wire ap_ST_fsm_state198_blk;
    wire ap_ST_fsm_state199_blk;
    wire ap_ST_fsm_state200_blk;
    wire ap_ST_fsm_state201_blk;
    wire ap_ST_fsm_state202_blk;
    wire ap_ST_fsm_state203_blk;
    reg ap_ST_fsm_state204_blk;
    wire ap_ST_fsm_state205_blk;
    wire ap_ST_fsm_state206_blk;
    reg ap_ST_fsm_state207_blk;
    wire ap_ST_fsm_state208_blk;
    reg ap_ST_fsm_state209_blk;
    wire ap_ST_fsm_state210_blk;
    wire ap_ST_fsm_state211_blk;
    wire ap_ST_fsm_state212_blk;
    wire ap_ST_fsm_state213_blk;
    wire ap_ST_fsm_state214_blk;
    wire ap_ST_fsm_state215_blk;
    reg ap_ST_fsm_state216_blk;
    reg ap_ST_fsm_state217_blk;
    wire ap_ST_fsm_state218_blk;
    wire ap_ST_fsm_state219_blk;
    wire ap_ST_fsm_state220_blk;
    wire ap_ST_fsm_state221_blk;
    wire ap_ST_fsm_state222_blk;
    wire ap_ST_fsm_state223_blk;
    wire ap_ST_fsm_state224_blk;
    wire ap_ST_fsm_state225_blk;
    wire ap_ST_fsm_state226_blk;
    wire ap_ST_fsm_state227_blk;
    wire ap_ST_fsm_state228_blk;
    wire ap_ST_fsm_state229_blk;
    wire ap_ST_fsm_state230_blk;
    wire ap_ST_fsm_state231_blk;
    wire ap_ST_fsm_state232_blk;
    wire ap_ST_fsm_state233_blk;
    wire ap_ST_fsm_state234_blk;
    wire ap_ST_fsm_state235_blk;
    wire ap_ST_fsm_state236_blk;
    wire ap_ST_fsm_state237_blk;
    wire ap_ST_fsm_state238_blk;
    wire ap_ST_fsm_state239_blk;
    wire ap_ST_fsm_state240_blk;
    wire ap_ST_fsm_state241_blk;
    wire ap_ST_fsm_state242_blk;
    wire ap_ST_fsm_state243_blk;
    wire ap_ST_fsm_state244_blk;
    wire ap_ST_fsm_state245_blk;
    wire ap_ST_fsm_state246_blk;
    wire ap_ST_fsm_state247_blk;
    wire ap_ST_fsm_state248_blk;
    wire ap_ST_fsm_state249_blk;
    wire ap_ST_fsm_state250_blk;
    wire ap_ST_fsm_state251_blk;
    wire ap_ST_fsm_state252_blk;
    wire ap_ST_fsm_state253_blk;
    wire ap_ST_fsm_state254_blk;
    wire ap_ST_fsm_state255_blk;
    wire ap_ST_fsm_state256_blk;
    wire ap_ST_fsm_state257_blk;
    wire ap_ST_fsm_state258_blk;
    wire ap_ST_fsm_state259_blk;
    wire ap_ST_fsm_state260_blk;
    wire ap_ST_fsm_state261_blk;
    wire ap_ST_fsm_state262_blk;
    wire ap_ST_fsm_state263_blk;
    wire ap_ST_fsm_state264_blk;
    wire ap_ST_fsm_state265_blk;
    wire ap_ST_fsm_state266_blk;
    wire ap_ST_fsm_state267_blk;
    wire ap_ST_fsm_state268_blk;
    wire ap_ST_fsm_state269_blk;
    wire ap_ST_fsm_state270_blk;
    wire ap_ST_fsm_state271_blk;
    wire ap_ST_fsm_state272_blk;
    wire ap_ST_fsm_state273_blk;
    wire ap_ST_fsm_state274_blk;
    wire ap_ST_fsm_state275_blk;
    reg ap_ST_fsm_state276_blk;
    wire ap_ST_fsm_state277_blk;
    reg ap_ST_fsm_state278_blk;
    wire ap_ST_fsm_state279_blk;
    wire ap_ST_fsm_state280_blk;
    wire ap_ST_fsm_state281_blk;
    wire ap_ST_fsm_state282_blk;
    wire ap_ST_fsm_state283_blk;
    wire ap_ST_fsm_state284_blk;
    wire ap_ST_fsm_state285_blk;
    wire ap_ST_fsm_state286_blk;
    wire ap_ST_fsm_state287_blk;
    wire ap_ST_fsm_state288_blk;
    wire ap_ST_fsm_state289_blk;
    wire ap_ST_fsm_state290_blk;
    wire ap_ST_fsm_state291_blk;
    wire ap_ST_fsm_state292_blk;
    wire ap_ST_fsm_state293_blk;
    wire ap_ST_fsm_state294_blk;
    wire ap_ST_fsm_state295_blk;
    wire ap_ST_fsm_state296_blk;
    wire ap_ST_fsm_state297_blk;
    wire ap_ST_fsm_state298_blk;
    wire ap_ST_fsm_state299_blk;
    wire ap_ST_fsm_state300_blk;
    wire ap_ST_fsm_state301_blk;
    wire ap_ST_fsm_state302_blk;
    wire ap_ST_fsm_state303_blk;
    wire ap_ST_fsm_state304_blk;
    wire ap_ST_fsm_state305_blk;
    wire ap_ST_fsm_state306_blk;
    wire ap_ST_fsm_state307_blk;
    wire ap_ST_fsm_state308_blk;
    wire ap_ST_fsm_state309_blk;
    wire ap_ST_fsm_state310_blk;
    wire ap_ST_fsm_state311_blk;
    wire ap_ST_fsm_state312_blk;
    wire ap_ST_fsm_state313_blk;
    wire ap_ST_fsm_state314_blk;
    wire ap_ST_fsm_state315_blk;
    wire ap_ST_fsm_state316_blk;
    wire ap_ST_fsm_state317_blk;
    wire ap_ST_fsm_state318_blk;
    wire ap_ST_fsm_state319_blk;
    wire ap_ST_fsm_state320_blk;
    wire ap_ST_fsm_state321_blk;
    wire ap_ST_fsm_state322_blk;
    wire ap_ST_fsm_state323_blk;
    wire ap_ST_fsm_state324_blk;
    wire ap_ST_fsm_state325_blk;
    wire ap_ST_fsm_state326_blk;
    wire ap_ST_fsm_state327_blk;
    wire ap_ST_fsm_state328_blk;
    wire ap_ST_fsm_state329_blk;
    wire ap_ST_fsm_state330_blk;
    wire ap_ST_fsm_state331_blk;
    wire ap_ST_fsm_state332_blk;
    wire ap_ST_fsm_state333_blk;
    wire ap_ST_fsm_state334_blk;
    wire ap_ST_fsm_state335_blk;
    wire ap_ST_fsm_state336_blk;
    wire ap_ST_fsm_state337_blk;
    reg ap_ST_fsm_state338_blk;
    wire ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 338'd1;
        #0 lfsr = 16'd44257;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg = 1'b0;
        #0 grp_detectCollNode_fu_1055_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg = 1'b0;
        #0 grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg = 1'b0;
        #0 numVertices_fu_520 = 32'd0;
    end

    main_planRRT_goal_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) goal_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(goal_address0),
        .ce0(goal_ce0),
        .q0(goal_q0)
    );

    main_planRRT_ang_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) ang_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(ang_address0),
        .ce0(ang_ce0),
        .we0(ang_we0),
        .d0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_d0),
        .q0(ang_q0)
    );

    main_planRRT_rrtVertices_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(6000),
        .AddressWidth(13)
    ) rrtVertices_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(rrtVertices_address0),
        .ce0(rrtVertices_ce0),
        .we0(rrtVertices_we0),
        .d0(rrtVertices_d0),
        .q0(rrtVertices_q0)
    );

    main_planRRT_ang_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) qRand_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(qRand_address0),
        .ce0(qRand_ce0),
        .we0(qRand_we0),
        .d0(qRand_d0),
        .q0(qRand_q0)
    );

    main_planRRT_ang_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) qNear_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(qNear_address0),
        .ce0(qNear_ce0),
        .we0(qNear_we0),
        .d0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_d0),
        .q0(qNear_q0)
    );

    main_planRRT_ang_RAM_AUTO_1R1W #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) qConnect_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(qConnect_address0),
        .ce0(qConnect_ce0),
        .we0(qConnect_we0),
        .d0(qConnect_d0),
        .q0(qConnect_q0)
    );

    main_planRRT_Pipeline_VITIS_LOOP_86_1 grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_ready),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_ce0),
        .rrtVertices_we0(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_we0),
        .rrtVertices_d0(grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_d0)
    );

    main_planRRT_Pipeline_VITIS_LOOP_152_1 grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_ready),
        .lfsr_load(lfsr),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_ce0),
        .qRand_we0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_we0),
        .qRand_d0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_d0),
        .or_i_i_i110_out(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out),
        .or_i_i_i110_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out_ap_vld),
        .shr6_i_i_i_phi_out(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out),
        .shr6_i_i_i_phi_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out_ap_vld),
        .grp_fu_1431_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din0),
        .grp_fu_1431_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din1),
        .grp_fu_1431_p_dout0(grp_fu_1431_p2),
        .grp_fu_1431_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_ce),
        .grp_fu_1436_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_din0),
        .grp_fu_1436_p_dout0(grp_fu_1436_p1),
        .grp_fu_1436_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_ce),
        .grp_fu_1439_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_din0),
        .grp_fu_1439_p_dout0(grp_fu_1439_p1),
        .grp_fu_1439_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_ce),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_110_4 grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_ready),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_ce0),
        .qRand_we0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_we0),
        .qRand_d0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_d0),
        .goal_address0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_address0),
        .goal_ce0(grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_ce0),
        .goal_q0(goal_q0)
    );

    main_planRRT_Pipeline_VITIS_LOOP_293_1 grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_ready),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_ce0),
        .qRand_q0(qRand_q0),
        .dist_out(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_dist_out),
        .dist_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_dist_out_ap_vld),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1 grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_ready),
        .minDist(reg_1470),
        .sub_ln296(sub_ln296_reg_2445),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_ce0),
        .qRand_q0(qRand_q0),
        .bestIdx_3_out(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out),
        .bestIdx_3_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out_ap_vld),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_ce),
        .grp_fu_1454_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din0),
        .grp_fu_1454_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din1),
        .grp_fu_1454_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_opcode),
        .grp_fu_1454_p_dout0(grp_fu_1454_p2),
        .grp_fu_1454_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_ce),
        .grp_fu_1462_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din0),
        .grp_fu_1462_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din1),
        .grp_fu_1462_p_dout0(grp_fu_1462_p2),
        .grp_fu_1462_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_114_5 grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_ready),
        .sub_ln114(sub_ln114_reg_2450),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .qNear_address0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_address0),
        .qNear_ce0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_ce0),
        .qNear_we0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_we0),
        .qNear_d0(grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_d0)
    );

    main_planRRT_Pipeline_VITIS_LOOP_293_18 grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_ready),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_ce0),
        .qRand_q0(qRand_q0),
        .qNear_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_address0),
        .qNear_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_ce0),
        .qNear_q0(qNear_q0),
        .dist_4_out(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_dist_4_out),
        .dist_4_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_dist_4_out_ap_vld),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_125_7 grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_ready),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_ce0),
        .qRand_q0(qRand_q0),
        .qConnect_address0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_address0),
        .qConnect_ce0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_ce0),
        .qConnect_we0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_we0),
        .qConnect_d0(grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_d0)
    );

    main_planRRT_Pipeline_VITIS_LOOP_121_6 grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_ready),
        .qNear_address0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_address0),
        .qNear_ce0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_ce0),
        .qNear_q0(qNear_q0),
        .qRand_address0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_address0),
        .qRand_ce0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_ce0),
        .qRand_q0(qRand_q0),
        .f(f_reg_2462),
        .qConnect_address0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_address0),
        .qConnect_ce0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_ce0),
        .qConnect_we0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_we0),
        .qConnect_d0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_d0),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_ce),
        .grp_fu_2537_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din0),
        .grp_fu_2537_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din1),
        .grp_fu_2537_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_opcode),
        .grp_fu_2537_p_dout0(grp_fu_2407_p_dout0),
        .grp_fu_2537_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_190_2 grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_ready),
        .qConnect_address0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_address0),
        .qConnect_ce0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_ce0),
        .qConnect_q0(qConnect_q0),
        .qNear_address0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_address0),
        .qNear_ce0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_ce0),
        .qNear_q0(qNear_q0),
        .s(s_reg_960),
        .ang_address0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_address0),
        .ang_ce0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_ce0),
        .ang_we0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_we0),
        .ang_d0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_d0),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_ce),
        .grp_fu_2537_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din0),
        .grp_fu_2537_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din1),
        .grp_fu_2537_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_opcode),
        .grp_fu_2537_p_dout0(grp_fu_2407_p_dout0),
        .grp_fu_2537_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_130_8 grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_ready),
        .sub_ln130(sub_ln130_reg_2431),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_ce0),
        .rrtVertices_we0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_we0),
        .rrtVertices_d0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_d0),
        .qConnect_address0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_address0),
        .qConnect_ce0(grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_ce0),
        .qConnect_q0(qConnect_q0)
    );

    main_detectCollNode grp_detectCollNode_fu_1055 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_detectCollNode_fu_1055_ap_start),
        .ap_done(grp_detectCollNode_fu_1055_ap_done),
        .ap_idle(grp_detectCollNode_fu_1055_ap_idle),
        .ap_ready(grp_detectCollNode_fu_1055_ap_ready),
        .this_env_0_0_0_address0(grp_detectCollNode_fu_1055_this_env_0_0_0_address0),
        .this_env_0_0_0_ce0(grp_detectCollNode_fu_1055_this_env_0_0_0_ce0),
        .this_env_0_0_0_q0(this_0_0_0_0_q0),
        .this_env_0_0_1_address0(grp_detectCollNode_fu_1055_this_env_0_0_1_address0),
        .this_env_0_0_1_ce0(grp_detectCollNode_fu_1055_this_env_0_0_1_ce0),
        .this_env_0_0_1_q0(this_0_0_0_1_q0),
        .this_env_0_0_2_address0(grp_detectCollNode_fu_1055_this_env_0_0_2_address0),
        .this_env_0_0_2_ce0(grp_detectCollNode_fu_1055_this_env_0_0_2_ce0),
        .this_env_0_0_2_q0(this_0_0_0_2_q0),
        .this_env_0_1_0_address0(grp_detectCollNode_fu_1055_this_env_0_1_0_address0),
        .this_env_0_1_0_ce0(grp_detectCollNode_fu_1055_this_env_0_1_0_ce0),
        .this_env_0_1_0_q0(this_0_0_1_0_q0),
        .this_env_0_1_1_address0(grp_detectCollNode_fu_1055_this_env_0_1_1_address0),
        .this_env_0_1_1_ce0(grp_detectCollNode_fu_1055_this_env_0_1_1_ce0),
        .this_env_0_1_1_q0(this_0_0_1_1_q0),
        .this_env_0_1_2_address0(grp_detectCollNode_fu_1055_this_env_0_1_2_address0),
        .this_env_0_1_2_ce0(grp_detectCollNode_fu_1055_this_env_0_1_2_ce0),
        .this_env_0_1_2_q0(this_0_0_1_2_q0),
        .this_env_0_2_0_address0(grp_detectCollNode_fu_1055_this_env_0_2_0_address0),
        .this_env_0_2_0_ce0(grp_detectCollNode_fu_1055_this_env_0_2_0_ce0),
        .this_env_0_2_0_q0(this_0_0_2_0_q0),
        .this_env_0_2_1_address0(grp_detectCollNode_fu_1055_this_env_0_2_1_address0),
        .this_env_0_2_1_ce0(grp_detectCollNode_fu_1055_this_env_0_2_1_ce0),
        .this_env_0_2_1_q0(this_0_0_2_1_q0),
        .this_env_0_2_2_address0(grp_detectCollNode_fu_1055_this_env_0_2_2_address0),
        .this_env_0_2_2_ce0(grp_detectCollNode_fu_1055_this_env_0_2_2_ce0),
        .this_env_0_2_2_q0(this_0_0_2_2_q0),
        .this_env_0_3_0_address0(grp_detectCollNode_fu_1055_this_env_0_3_0_address0),
        .this_env_0_3_0_ce0(grp_detectCollNode_fu_1055_this_env_0_3_0_ce0),
        .this_env_0_3_0_q0(this_0_0_3_0_q0),
        .this_env_0_3_1_address0(grp_detectCollNode_fu_1055_this_env_0_3_1_address0),
        .this_env_0_3_1_ce0(grp_detectCollNode_fu_1055_this_env_0_3_1_ce0),
        .this_env_0_3_1_q0(this_0_0_3_1_q0),
        .this_env_0_3_2_address0(grp_detectCollNode_fu_1055_this_env_0_3_2_address0),
        .this_env_0_3_2_ce0(grp_detectCollNode_fu_1055_this_env_0_3_2_ce0),
        .this_env_0_3_2_q0(this_0_0_3_2_q0),
        .this_env_0_4_0_address0(grp_detectCollNode_fu_1055_this_env_0_4_0_address0),
        .this_env_0_4_0_ce0(grp_detectCollNode_fu_1055_this_env_0_4_0_ce0),
        .this_env_0_4_0_q0(this_0_0_4_0_q0),
        .this_env_0_4_1_address0(grp_detectCollNode_fu_1055_this_env_0_4_1_address0),
        .this_env_0_4_1_ce0(grp_detectCollNode_fu_1055_this_env_0_4_1_ce0),
        .this_env_0_4_1_q0(this_0_0_4_1_q0),
        .this_env_0_4_2_address0(grp_detectCollNode_fu_1055_this_env_0_4_2_address0),
        .this_env_0_4_2_ce0(grp_detectCollNode_fu_1055_this_env_0_4_2_ce0),
        .this_env_0_4_2_q0(this_0_0_4_2_q0),
        .this_env_0_5_0_address0(grp_detectCollNode_fu_1055_this_env_0_5_0_address0),
        .this_env_0_5_0_ce0(grp_detectCollNode_fu_1055_this_env_0_5_0_ce0),
        .this_env_0_5_0_q0(this_0_0_5_0_q0),
        .this_env_0_5_1_address0(grp_detectCollNode_fu_1055_this_env_0_5_1_address0),
        .this_env_0_5_1_ce0(grp_detectCollNode_fu_1055_this_env_0_5_1_ce0),
        .this_env_0_5_1_q0(this_0_0_5_1_q0),
        .this_env_0_5_2_address0(grp_detectCollNode_fu_1055_this_env_0_5_2_address0),
        .this_env_0_5_2_ce0(grp_detectCollNode_fu_1055_this_env_0_5_2_ce0),
        .this_env_0_5_2_q0(this_0_0_5_2_q0),
        .this_env_0_6_0_address0(grp_detectCollNode_fu_1055_this_env_0_6_0_address0),
        .this_env_0_6_0_ce0(grp_detectCollNode_fu_1055_this_env_0_6_0_ce0),
        .this_env_0_6_0_q0(this_0_0_6_0_q0),
        .this_env_0_6_1_address0(grp_detectCollNode_fu_1055_this_env_0_6_1_address0),
        .this_env_0_6_1_ce0(grp_detectCollNode_fu_1055_this_env_0_6_1_ce0),
        .this_env_0_6_1_q0(this_0_0_6_1_q0),
        .this_env_0_6_2_address0(grp_detectCollNode_fu_1055_this_env_0_6_2_address0),
        .this_env_0_6_2_ce0(grp_detectCollNode_fu_1055_this_env_0_6_2_ce0),
        .this_env_0_6_2_q0(this_0_0_6_2_q0),
        .this_env_0_7_0_address0(grp_detectCollNode_fu_1055_this_env_0_7_0_address0),
        .this_env_0_7_0_ce0(grp_detectCollNode_fu_1055_this_env_0_7_0_ce0),
        .this_env_0_7_0_q0(this_0_0_7_0_q0),
        .this_env_0_7_1_address0(grp_detectCollNode_fu_1055_this_env_0_7_1_address0),
        .this_env_0_7_1_ce0(grp_detectCollNode_fu_1055_this_env_0_7_1_ce0),
        .this_env_0_7_1_q0(this_0_0_7_1_q0),
        .this_env_0_7_2_address0(grp_detectCollNode_fu_1055_this_env_0_7_2_address0),
        .this_env_0_7_2_ce0(grp_detectCollNode_fu_1055_this_env_0_7_2_ce0),
        .this_env_0_7_2_q0(this_0_0_7_2_q0),
        .this_env_0_8_0_address0(grp_detectCollNode_fu_1055_this_env_0_8_0_address0),
        .this_env_0_8_0_ce0(grp_detectCollNode_fu_1055_this_env_0_8_0_ce0),
        .this_env_0_8_0_q0(this_0_0_8_0_q0),
        .this_env_0_8_1_address0(grp_detectCollNode_fu_1055_this_env_0_8_1_address0),
        .this_env_0_8_1_ce0(grp_detectCollNode_fu_1055_this_env_0_8_1_ce0),
        .this_env_0_8_1_q0(this_0_0_8_1_q0),
        .this_env_0_8_2_address0(grp_detectCollNode_fu_1055_this_env_0_8_2_address0),
        .this_env_0_8_2_ce0(grp_detectCollNode_fu_1055_this_env_0_8_2_ce0),
        .this_env_0_8_2_q0(this_0_0_8_2_q0),
        .this_env_1_address0(grp_detectCollNode_fu_1055_this_env_1_address0),
        .this_env_1_ce0(grp_detectCollNode_fu_1055_this_env_1_ce0),
        .this_env_1_q0(this_0_1_q0),
        .this_env_1_address1(grp_detectCollNode_fu_1055_this_env_1_address1),
        .this_env_1_ce1(grp_detectCollNode_fu_1055_this_env_1_ce1),
        .this_env_1_q1(this_0_1_q1),
        .this_TLink_0_0_address0(grp_detectCollNode_fu_1055_this_TLink_0_0_address0),
        .this_TLink_0_0_ce0(grp_detectCollNode_fu_1055_this_TLink_0_0_ce0),
        .this_TLink_0_0_q0(this_4_0_0_q0),
        .this_TLink_0_1_address0(grp_detectCollNode_fu_1055_this_TLink_0_1_address0),
        .this_TLink_0_1_ce0(grp_detectCollNode_fu_1055_this_TLink_0_1_ce0),
        .this_TLink_0_1_q0(this_4_0_1_q0),
        .this_TLink_0_2_address0(grp_detectCollNode_fu_1055_this_TLink_0_2_address0),
        .this_TLink_0_2_ce0(grp_detectCollNode_fu_1055_this_TLink_0_2_ce0),
        .this_TLink_0_2_q0(this_4_0_2_q0),
        .this_TLink_0_3_address0(grp_detectCollNode_fu_1055_this_TLink_0_3_address0),
        .this_TLink_0_3_ce0(grp_detectCollNode_fu_1055_this_TLink_0_3_ce0),
        .this_TLink_0_3_q0(this_4_0_3_q0),
        .this_TLink_1_0_address0(grp_detectCollNode_fu_1055_this_TLink_1_0_address0),
        .this_TLink_1_0_ce0(grp_detectCollNode_fu_1055_this_TLink_1_0_ce0),
        .this_TLink_1_0_q0(this_4_1_0_q0),
        .this_TLink_1_1_address0(grp_detectCollNode_fu_1055_this_TLink_1_1_address0),
        .this_TLink_1_1_ce0(grp_detectCollNode_fu_1055_this_TLink_1_1_ce0),
        .this_TLink_1_1_q0(this_4_1_1_q0),
        .this_TLink_1_2_address0(grp_detectCollNode_fu_1055_this_TLink_1_2_address0),
        .this_TLink_1_2_ce0(grp_detectCollNode_fu_1055_this_TLink_1_2_ce0),
        .this_TLink_1_2_q0(this_4_1_2_q0),
        .this_TLink_1_3_address0(grp_detectCollNode_fu_1055_this_TLink_1_3_address0),
        .this_TLink_1_3_ce0(grp_detectCollNode_fu_1055_this_TLink_1_3_ce0),
        .this_TLink_1_3_q0(this_4_1_3_q0),
        .this_TLink_2_0_address0(grp_detectCollNode_fu_1055_this_TLink_2_0_address0),
        .this_TLink_2_0_ce0(grp_detectCollNode_fu_1055_this_TLink_2_0_ce0),
        .this_TLink_2_0_q0(this_4_2_0_q0),
        .this_TLink_2_1_address0(grp_detectCollNode_fu_1055_this_TLink_2_1_address0),
        .this_TLink_2_1_ce0(grp_detectCollNode_fu_1055_this_TLink_2_1_ce0),
        .this_TLink_2_1_q0(this_4_2_1_q0),
        .this_TLink_2_2_address0(grp_detectCollNode_fu_1055_this_TLink_2_2_address0),
        .this_TLink_2_2_ce0(grp_detectCollNode_fu_1055_this_TLink_2_2_ce0),
        .this_TLink_2_2_q0(this_4_2_2_q0),
        .this_TLink_2_3_address0(grp_detectCollNode_fu_1055_this_TLink_2_3_address0),
        .this_TLink_2_3_ce0(grp_detectCollNode_fu_1055_this_TLink_2_3_ce0),
        .this_TLink_2_3_q0(this_4_2_3_q0),
        .this_TLink_3_0_address0(grp_detectCollNode_fu_1055_this_TLink_3_0_address0),
        .this_TLink_3_0_ce0(grp_detectCollNode_fu_1055_this_TLink_3_0_ce0),
        .this_TLink_3_0_q0(this_4_3_0_q0),
        .this_TLink_3_1_address0(grp_detectCollNode_fu_1055_this_TLink_3_1_address0),
        .this_TLink_3_1_ce0(grp_detectCollNode_fu_1055_this_TLink_3_1_ce0),
        .this_TLink_3_1_q0(this_4_3_1_q0),
        .this_TLink_3_2_address0(grp_detectCollNode_fu_1055_this_TLink_3_2_address0),
        .this_TLink_3_2_ce0(grp_detectCollNode_fu_1055_this_TLink_3_2_ce0),
        .this_TLink_3_2_q0(this_4_3_2_q0),
        .this_TLink_3_3_address0(grp_detectCollNode_fu_1055_this_TLink_3_3_address0),
        .this_TLink_3_3_ce0(grp_detectCollNode_fu_1055_this_TLink_3_3_ce0),
        .this_TLink_3_3_q0(this_4_3_3_q0),
        .this_TJoint_0_0_address0(grp_detectCollNode_fu_1055_this_TJoint_0_0_address0),
        .this_TJoint_0_0_ce0(grp_detectCollNode_fu_1055_this_TJoint_0_0_ce0),
        .this_TJoint_0_0_we0(grp_detectCollNode_fu_1055_this_TJoint_0_0_we0),
        .this_TJoint_0_0_d0(grp_detectCollNode_fu_1055_this_TJoint_0_0_d0),
        .this_TJoint_0_0_q0(this_5_0_0_q0),
        .this_TJoint_0_1_address0(grp_detectCollNode_fu_1055_this_TJoint_0_1_address0),
        .this_TJoint_0_1_ce0(grp_detectCollNode_fu_1055_this_TJoint_0_1_ce0),
        .this_TJoint_0_1_we0(grp_detectCollNode_fu_1055_this_TJoint_0_1_we0),
        .this_TJoint_0_1_d0(grp_detectCollNode_fu_1055_this_TJoint_0_1_d0),
        .this_TJoint_0_1_q0(this_5_0_1_q0),
        .this_TJoint_0_2_address0(grp_detectCollNode_fu_1055_this_TJoint_0_2_address0),
        .this_TJoint_0_2_ce0(grp_detectCollNode_fu_1055_this_TJoint_0_2_ce0),
        .this_TJoint_0_2_we0(grp_detectCollNode_fu_1055_this_TJoint_0_2_we0),
        .this_TJoint_0_2_d0(grp_detectCollNode_fu_1055_this_TJoint_0_2_d0),
        .this_TJoint_0_2_q0(this_5_0_2_q0),
        .this_TJoint_0_3_address0(grp_detectCollNode_fu_1055_this_TJoint_0_3_address0),
        .this_TJoint_0_3_ce0(grp_detectCollNode_fu_1055_this_TJoint_0_3_ce0),
        .this_TJoint_0_3_we0(grp_detectCollNode_fu_1055_this_TJoint_0_3_we0),
        .this_TJoint_0_3_d0(grp_detectCollNode_fu_1055_this_TJoint_0_3_d0),
        .this_TJoint_0_3_q0(this_5_0_3_q0),
        .this_TJoint_1_0_address0(grp_detectCollNode_fu_1055_this_TJoint_1_0_address0),
        .this_TJoint_1_0_ce0(grp_detectCollNode_fu_1055_this_TJoint_1_0_ce0),
        .this_TJoint_1_0_we0(grp_detectCollNode_fu_1055_this_TJoint_1_0_we0),
        .this_TJoint_1_0_d0(grp_detectCollNode_fu_1055_this_TJoint_1_0_d0),
        .this_TJoint_1_0_q0(this_5_1_0_q0),
        .this_TJoint_1_1_address0(grp_detectCollNode_fu_1055_this_TJoint_1_1_address0),
        .this_TJoint_1_1_ce0(grp_detectCollNode_fu_1055_this_TJoint_1_1_ce0),
        .this_TJoint_1_1_we0(grp_detectCollNode_fu_1055_this_TJoint_1_1_we0),
        .this_TJoint_1_1_d0(grp_detectCollNode_fu_1055_this_TJoint_1_1_d0),
        .this_TJoint_1_1_q0(this_5_1_1_q0),
        .this_TJoint_1_2_address0(grp_detectCollNode_fu_1055_this_TJoint_1_2_address0),
        .this_TJoint_1_2_ce0(grp_detectCollNode_fu_1055_this_TJoint_1_2_ce0),
        .this_TJoint_1_2_we0(grp_detectCollNode_fu_1055_this_TJoint_1_2_we0),
        .this_TJoint_1_2_d0(grp_detectCollNode_fu_1055_this_TJoint_1_2_d0),
        .this_TJoint_1_2_q0(this_5_1_2_q0),
        .this_TJoint_1_3_address0(grp_detectCollNode_fu_1055_this_TJoint_1_3_address0),
        .this_TJoint_1_3_ce0(grp_detectCollNode_fu_1055_this_TJoint_1_3_ce0),
        .this_TJoint_1_3_we0(grp_detectCollNode_fu_1055_this_TJoint_1_3_we0),
        .this_TJoint_1_3_d0(grp_detectCollNode_fu_1055_this_TJoint_1_3_d0),
        .this_TJoint_1_3_q0(this_5_1_3_q0),
        .this_TJoint_2_0_address0(grp_detectCollNode_fu_1055_this_TJoint_2_0_address0),
        .this_TJoint_2_0_ce0(grp_detectCollNode_fu_1055_this_TJoint_2_0_ce0),
        .this_TJoint_2_0_we0(grp_detectCollNode_fu_1055_this_TJoint_2_0_we0),
        .this_TJoint_2_0_d0(grp_detectCollNode_fu_1055_this_TJoint_2_0_d0),
        .this_TJoint_2_0_q0(this_5_2_0_q0),
        .this_TJoint_2_1_address0(grp_detectCollNode_fu_1055_this_TJoint_2_1_address0),
        .this_TJoint_2_1_ce0(grp_detectCollNode_fu_1055_this_TJoint_2_1_ce0),
        .this_TJoint_2_1_we0(grp_detectCollNode_fu_1055_this_TJoint_2_1_we0),
        .this_TJoint_2_1_d0(grp_detectCollNode_fu_1055_this_TJoint_2_1_d0),
        .this_TJoint_2_1_q0(this_5_2_1_q0),
        .this_TJoint_2_2_address0(grp_detectCollNode_fu_1055_this_TJoint_2_2_address0),
        .this_TJoint_2_2_ce0(grp_detectCollNode_fu_1055_this_TJoint_2_2_ce0),
        .this_TJoint_2_2_we0(grp_detectCollNode_fu_1055_this_TJoint_2_2_we0),
        .this_TJoint_2_2_d0(grp_detectCollNode_fu_1055_this_TJoint_2_2_d0),
        .this_TJoint_2_2_q0(this_5_2_2_q0),
        .this_TJoint_2_3_address0(grp_detectCollNode_fu_1055_this_TJoint_2_3_address0),
        .this_TJoint_2_3_ce0(grp_detectCollNode_fu_1055_this_TJoint_2_3_ce0),
        .this_TJoint_2_3_we0(grp_detectCollNode_fu_1055_this_TJoint_2_3_we0),
        .this_TJoint_2_3_d0(grp_detectCollNode_fu_1055_this_TJoint_2_3_d0),
        .this_TJoint_2_3_q0(this_5_2_3_q0),
        .this_TJoint_3_0_address0(grp_detectCollNode_fu_1055_this_TJoint_3_0_address0),
        .this_TJoint_3_0_ce0(grp_detectCollNode_fu_1055_this_TJoint_3_0_ce0),
        .this_TJoint_3_0_we0(grp_detectCollNode_fu_1055_this_TJoint_3_0_we0),
        .this_TJoint_3_0_d0(grp_detectCollNode_fu_1055_this_TJoint_3_0_d0),
        .this_TJoint_3_0_q0(this_5_3_0_q0),
        .this_TJoint_3_1_address0(grp_detectCollNode_fu_1055_this_TJoint_3_1_address0),
        .this_TJoint_3_1_ce0(grp_detectCollNode_fu_1055_this_TJoint_3_1_ce0),
        .this_TJoint_3_1_we0(grp_detectCollNode_fu_1055_this_TJoint_3_1_we0),
        .this_TJoint_3_1_d0(grp_detectCollNode_fu_1055_this_TJoint_3_1_d0),
        .this_TJoint_3_1_q0(this_5_3_1_q0),
        .this_TJoint_3_2_address0(grp_detectCollNode_fu_1055_this_TJoint_3_2_address0),
        .this_TJoint_3_2_ce0(grp_detectCollNode_fu_1055_this_TJoint_3_2_ce0),
        .this_TJoint_3_2_we0(grp_detectCollNode_fu_1055_this_TJoint_3_2_we0),
        .this_TJoint_3_2_d0(grp_detectCollNode_fu_1055_this_TJoint_3_2_d0),
        .this_TJoint_3_2_q0(this_5_3_2_q0),
        .this_TJoint_3_3_address0(grp_detectCollNode_fu_1055_this_TJoint_3_3_address0),
        .this_TJoint_3_3_ce0(grp_detectCollNode_fu_1055_this_TJoint_3_3_ce0),
        .this_TJoint_3_3_we0(grp_detectCollNode_fu_1055_this_TJoint_3_3_we0),
        .this_TJoint_3_3_d0(grp_detectCollNode_fu_1055_this_TJoint_3_3_d0),
        .this_TJoint_3_3_q0(this_5_3_3_q0),
        .this_TCurr_0_0_address0(grp_detectCollNode_fu_1055_this_TCurr_0_0_address0),
        .this_TCurr_0_0_ce0(grp_detectCollNode_fu_1055_this_TCurr_0_0_ce0),
        .this_TCurr_0_0_we0(grp_detectCollNode_fu_1055_this_TCurr_0_0_we0),
        .this_TCurr_0_0_d0(grp_detectCollNode_fu_1055_this_TCurr_0_0_d0),
        .this_TCurr_0_0_q0(this_6_0_0_q0),
        .this_TCurr_0_1_address0(grp_detectCollNode_fu_1055_this_TCurr_0_1_address0),
        .this_TCurr_0_1_ce0(grp_detectCollNode_fu_1055_this_TCurr_0_1_ce0),
        .this_TCurr_0_1_we0(grp_detectCollNode_fu_1055_this_TCurr_0_1_we0),
        .this_TCurr_0_1_d0(grp_detectCollNode_fu_1055_this_TCurr_0_1_d0),
        .this_TCurr_0_1_q0(this_6_0_1_q0),
        .this_TCurr_0_2_address0(grp_detectCollNode_fu_1055_this_TCurr_0_2_address0),
        .this_TCurr_0_2_ce0(grp_detectCollNode_fu_1055_this_TCurr_0_2_ce0),
        .this_TCurr_0_2_we0(grp_detectCollNode_fu_1055_this_TCurr_0_2_we0),
        .this_TCurr_0_2_d0(grp_detectCollNode_fu_1055_this_TCurr_0_2_d0),
        .this_TCurr_0_2_q0(this_6_0_2_q0),
        .this_TCurr_0_3_address0(grp_detectCollNode_fu_1055_this_TCurr_0_3_address0),
        .this_TCurr_0_3_ce0(grp_detectCollNode_fu_1055_this_TCurr_0_3_ce0),
        .this_TCurr_0_3_we0(grp_detectCollNode_fu_1055_this_TCurr_0_3_we0),
        .this_TCurr_0_3_d0(grp_detectCollNode_fu_1055_this_TCurr_0_3_d0),
        .this_TCurr_0_3_q0(this_6_0_3_q0),
        .this_TCurr_1_0_address0(grp_detectCollNode_fu_1055_this_TCurr_1_0_address0),
        .this_TCurr_1_0_ce0(grp_detectCollNode_fu_1055_this_TCurr_1_0_ce0),
        .this_TCurr_1_0_we0(grp_detectCollNode_fu_1055_this_TCurr_1_0_we0),
        .this_TCurr_1_0_d0(grp_detectCollNode_fu_1055_this_TCurr_1_0_d0),
        .this_TCurr_1_0_q0(this_6_1_0_q0),
        .this_TCurr_1_1_address0(grp_detectCollNode_fu_1055_this_TCurr_1_1_address0),
        .this_TCurr_1_1_ce0(grp_detectCollNode_fu_1055_this_TCurr_1_1_ce0),
        .this_TCurr_1_1_we0(grp_detectCollNode_fu_1055_this_TCurr_1_1_we0),
        .this_TCurr_1_1_d0(grp_detectCollNode_fu_1055_this_TCurr_1_1_d0),
        .this_TCurr_1_1_q0(this_6_1_1_q0),
        .this_TCurr_1_2_address0(grp_detectCollNode_fu_1055_this_TCurr_1_2_address0),
        .this_TCurr_1_2_ce0(grp_detectCollNode_fu_1055_this_TCurr_1_2_ce0),
        .this_TCurr_1_2_we0(grp_detectCollNode_fu_1055_this_TCurr_1_2_we0),
        .this_TCurr_1_2_d0(grp_detectCollNode_fu_1055_this_TCurr_1_2_d0),
        .this_TCurr_1_2_q0(this_6_1_2_q0),
        .this_TCurr_1_3_address0(grp_detectCollNode_fu_1055_this_TCurr_1_3_address0),
        .this_TCurr_1_3_ce0(grp_detectCollNode_fu_1055_this_TCurr_1_3_ce0),
        .this_TCurr_1_3_we0(grp_detectCollNode_fu_1055_this_TCurr_1_3_we0),
        .this_TCurr_1_3_d0(grp_detectCollNode_fu_1055_this_TCurr_1_3_d0),
        .this_TCurr_1_3_q0(this_6_1_3_q0),
        .this_TCurr_2_0_address0(grp_detectCollNode_fu_1055_this_TCurr_2_0_address0),
        .this_TCurr_2_0_ce0(grp_detectCollNode_fu_1055_this_TCurr_2_0_ce0),
        .this_TCurr_2_0_we0(grp_detectCollNode_fu_1055_this_TCurr_2_0_we0),
        .this_TCurr_2_0_d0(grp_detectCollNode_fu_1055_this_TCurr_2_0_d0),
        .this_TCurr_2_0_q0(this_6_2_0_q0),
        .this_TCurr_2_1_address0(grp_detectCollNode_fu_1055_this_TCurr_2_1_address0),
        .this_TCurr_2_1_ce0(grp_detectCollNode_fu_1055_this_TCurr_2_1_ce0),
        .this_TCurr_2_1_we0(grp_detectCollNode_fu_1055_this_TCurr_2_1_we0),
        .this_TCurr_2_1_d0(grp_detectCollNode_fu_1055_this_TCurr_2_1_d0),
        .this_TCurr_2_1_q0(this_6_2_1_q0),
        .this_TCurr_2_2_address0(grp_detectCollNode_fu_1055_this_TCurr_2_2_address0),
        .this_TCurr_2_2_ce0(grp_detectCollNode_fu_1055_this_TCurr_2_2_ce0),
        .this_TCurr_2_2_we0(grp_detectCollNode_fu_1055_this_TCurr_2_2_we0),
        .this_TCurr_2_2_d0(grp_detectCollNode_fu_1055_this_TCurr_2_2_d0),
        .this_TCurr_2_2_q0(this_6_2_2_q0),
        .this_TCurr_2_3_address0(grp_detectCollNode_fu_1055_this_TCurr_2_3_address0),
        .this_TCurr_2_3_ce0(grp_detectCollNode_fu_1055_this_TCurr_2_3_ce0),
        .this_TCurr_2_3_we0(grp_detectCollNode_fu_1055_this_TCurr_2_3_we0),
        .this_TCurr_2_3_d0(grp_detectCollNode_fu_1055_this_TCurr_2_3_d0),
        .this_TCurr_2_3_q0(this_6_2_3_q0),
        .this_TCurr_3_0_address0(grp_detectCollNode_fu_1055_this_TCurr_3_0_address0),
        .this_TCurr_3_0_ce0(grp_detectCollNode_fu_1055_this_TCurr_3_0_ce0),
        .this_TCurr_3_0_we0(grp_detectCollNode_fu_1055_this_TCurr_3_0_we0),
        .this_TCurr_3_0_d0(grp_detectCollNode_fu_1055_this_TCurr_3_0_d0),
        .this_TCurr_3_0_q0(this_6_3_0_q0),
        .this_TCurr_3_1_address0(grp_detectCollNode_fu_1055_this_TCurr_3_1_address0),
        .this_TCurr_3_1_ce0(grp_detectCollNode_fu_1055_this_TCurr_3_1_ce0),
        .this_TCurr_3_1_we0(grp_detectCollNode_fu_1055_this_TCurr_3_1_we0),
        .this_TCurr_3_1_d0(grp_detectCollNode_fu_1055_this_TCurr_3_1_d0),
        .this_TCurr_3_1_q0(this_6_3_1_q0),
        .this_TCurr_3_2_address0(grp_detectCollNode_fu_1055_this_TCurr_3_2_address0),
        .this_TCurr_3_2_ce0(grp_detectCollNode_fu_1055_this_TCurr_3_2_ce0),
        .this_TCurr_3_2_we0(grp_detectCollNode_fu_1055_this_TCurr_3_2_we0),
        .this_TCurr_3_2_d0(grp_detectCollNode_fu_1055_this_TCurr_3_2_d0),
        .this_TCurr_3_2_q0(this_6_3_2_q0),
        .this_TCurr_3_3_address0(grp_detectCollNode_fu_1055_this_TCurr_3_3_address0),
        .this_TCurr_3_3_ce0(grp_detectCollNode_fu_1055_this_TCurr_3_3_ce0),
        .this_TCurr_3_3_we0(grp_detectCollNode_fu_1055_this_TCurr_3_3_we0),
        .this_TCurr_3_3_d0(grp_detectCollNode_fu_1055_this_TCurr_3_3_d0),
        .this_TCurr_3_3_q0(this_6_3_3_q0),
        .this_q_address0(grp_detectCollNode_fu_1055_this_q_address0),
        .this_q_ce0(grp_detectCollNode_fu_1055_this_q_ce0),
        .this_q_we0(grp_detectCollNode_fu_1055_this_q_we0),
        .this_q_d0(grp_detectCollNode_fu_1055_this_q_d0),
        .this_q_q0(this_7_q0),
        .p_read(p_read),
        .p_read1(p_read1),
        .p_read2(p_read2),
        .p_read3(p_read3),
        .p_read4(p_read4),
        .p_read5(p_read5),
        .p_read6(p_read6),
        .p_read7(p_read7),
        .p_read8(p_read8),
        .p_read9(p_read9),
        .p_read10(p_read10),
        .p_read11(p_read11),
        .p_read12(p_read12),
        .p_read13(p_read13),
        .p_read14(p_read14),
        .p_read15(p_read15),
        .p_read16(p_read16),
        .p_read17(p_read17),
        .p_read18(p_read18),
        .p_read19(p_read19),
        .p_read20(p_read20),
        .p_read21(p_read21),
        .p_read22(p_read22),
        .p_read23(p_read23),
        .p_read24(p_read24),
        .p_read25(p_read25),
        .p_read26(p_read26),
        .p_read27(p_read27),
        .p_read28(p_read28),
        .p_read29(p_read29),
        .p_read30(p_read30),
        .p_read31(p_read31),
        .p_read32(p_read32),
        .p_read33(p_read33),
        .p_read34(p_read34),
        .p_read35(p_read35),
        .p_read36(p_read36),
        .p_read37(p_read37),
        .p_read38(p_read38),
        .p_read39(p_read39),
        .p_read40(p_read40),
        .p_read41(p_read41),
        .p_read42(p_read42),
        .p_read43(p_read43),
        .p_read44(p_read44),
        .p_read45(p_read45),
        .p_read46(p_read46),
        .p_read47(p_read47),
        .p_read48(p_read48),
        .p_read49(p_read49),
        .p_read50(p_read50),
        .p_read51(p_read51),
        .p_read52(p_read52),
        .p_read53(p_read53),
        .p_read54(p_read54),
        .p_read55(p_read55),
        .p_read56(p_read56),
        .p_read57(p_read57),
        .p_read58(p_read58),
        .p_read59(p_read59),
        .p_read60(p_read60),
        .p_read61(p_read61),
        .p_read62(p_read62),
        .p_read63(p_read63),
        .this_cPoints_address0(grp_detectCollNode_fu_1055_this_cPoints_address0),
        .this_cPoints_ce0(grp_detectCollNode_fu_1055_this_cPoints_ce0),
        .this_cPoints_we0(grp_detectCollNode_fu_1055_this_cPoints_we0),
        .this_cPoints_d0(grp_detectCollNode_fu_1055_this_cPoints_d0),
        .this_cPoints_q0(this_15_q0),
        .this_cPoints_address1(grp_detectCollNode_fu_1055_this_cPoints_address1),
        .this_cPoints_ce1(grp_detectCollNode_fu_1055_this_cPoints_ce1),
        .this_cPoints_we1(grp_detectCollNode_fu_1055_this_cPoints_we1),
        .this_cPoints_d1(grp_detectCollNode_fu_1055_this_cPoints_d1),
        .this_cPoints_q1(this_15_q1),
        .this_cAxes_address0(grp_detectCollNode_fu_1055_this_cAxes_address0),
        .this_cAxes_ce0(grp_detectCollNode_fu_1055_this_cAxes_ce0),
        .this_cAxes_we0(grp_detectCollNode_fu_1055_this_cAxes_we0),
        .this_cAxes_d0(grp_detectCollNode_fu_1055_this_cAxes_d0),
        .this_cAxes_q0(this_16_q0),
        .this_cAxes_address1(grp_detectCollNode_fu_1055_this_cAxes_address1),
        .this_cAxes_ce1(grp_detectCollNode_fu_1055_this_cAxes_ce1),
        .this_cAxes_q1(this_16_q1),
        .ang_address0(grp_detectCollNode_fu_1055_ang_address0),
        .ang_ce0(grp_detectCollNode_fu_1055_ang_ce0),
        .ang_q0(ang_q0),
        .l_TColl_0_0_0_constprop_i(l_TColl_0_0_0_constprop_i),
        .l_TColl_0_0_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o),
        .l_TColl_0_0_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o_ap_vld),
        .l_TColl_0_0_1_constprop_i(l_TColl_0_0_1_constprop_i),
        .l_TColl_0_0_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o),
        .l_TColl_0_0_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o_ap_vld),
        .l_TColl_0_0_2_constprop_i(l_TColl_0_0_2_constprop_i),
        .l_TColl_0_0_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o),
        .l_TColl_0_0_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o_ap_vld),
        .l_TColl_0_0_3_constprop_i(l_TColl_0_0_3_constprop_i),
        .l_TColl_0_0_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o),
        .l_TColl_0_0_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o_ap_vld),
        .l_TColl_1_0_0_constprop_i(l_TColl_1_0_0_constprop_i),
        .l_TColl_1_0_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o),
        .l_TColl_1_0_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o_ap_vld),
        .l_TColl_1_0_1_constprop_i(l_TColl_1_0_1_constprop_i),
        .l_TColl_1_0_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o),
        .l_TColl_1_0_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o_ap_vld),
        .l_TColl_1_0_2_constprop_i(l_TColl_1_0_2_constprop_i),
        .l_TColl_1_0_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o),
        .l_TColl_1_0_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o_ap_vld),
        .l_TColl_1_0_3_constprop_i(l_TColl_1_0_3_constprop_i),
        .l_TColl_1_0_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o),
        .l_TColl_1_0_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o_ap_vld),
        .l_TColl_2_0_0_constprop_i(l_TColl_2_0_0_constprop_i),
        .l_TColl_2_0_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o),
        .l_TColl_2_0_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o_ap_vld),
        .l_TColl_2_0_1_constprop_i(l_TColl_2_0_1_constprop_i),
        .l_TColl_2_0_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o),
        .l_TColl_2_0_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o_ap_vld),
        .l_TColl_2_0_2_constprop_i(l_TColl_2_0_2_constprop_i),
        .l_TColl_2_0_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o),
        .l_TColl_2_0_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o_ap_vld),
        .l_TColl_2_0_3_constprop_i(l_TColl_2_0_3_constprop_i),
        .l_TColl_2_0_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o),
        .l_TColl_2_0_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o_ap_vld),
        .l_TColl_0_1_0_constprop_i(l_TColl_0_1_0_constprop_i),
        .l_TColl_0_1_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o),
        .l_TColl_0_1_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o_ap_vld),
        .l_TColl_0_1_1_constprop_i(l_TColl_0_1_1_constprop_i),
        .l_TColl_0_1_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o),
        .l_TColl_0_1_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o_ap_vld),
        .l_TColl_0_1_2_constprop_i(l_TColl_0_1_2_constprop_i),
        .l_TColl_0_1_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o),
        .l_TColl_0_1_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o_ap_vld),
        .l_TColl_0_1_3_constprop_i(l_TColl_0_1_3_constprop_i),
        .l_TColl_0_1_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o),
        .l_TColl_0_1_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o_ap_vld),
        .l_TColl_1_1_0_constprop_i(l_TColl_1_1_0_constprop_i),
        .l_TColl_1_1_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o),
        .l_TColl_1_1_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o_ap_vld),
        .l_TColl_1_1_1_constprop_i(l_TColl_1_1_1_constprop_i),
        .l_TColl_1_1_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o),
        .l_TColl_1_1_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o_ap_vld),
        .l_TColl_1_1_2_constprop_i(l_TColl_1_1_2_constprop_i),
        .l_TColl_1_1_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o),
        .l_TColl_1_1_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o_ap_vld),
        .l_TColl_1_1_3_constprop_i(l_TColl_1_1_3_constprop_i),
        .l_TColl_1_1_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o),
        .l_TColl_1_1_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o_ap_vld),
        .l_TColl_2_1_0_constprop_i(l_TColl_2_1_0_constprop_i),
        .l_TColl_2_1_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o),
        .l_TColl_2_1_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o_ap_vld),
        .l_TColl_2_1_1_constprop_i(l_TColl_2_1_1_constprop_i),
        .l_TColl_2_1_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o),
        .l_TColl_2_1_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o_ap_vld),
        .l_TColl_2_1_2_constprop_i(l_TColl_2_1_2_constprop_i),
        .l_TColl_2_1_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o),
        .l_TColl_2_1_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o_ap_vld),
        .l_TColl_2_1_3_constprop_i(l_TColl_2_1_3_constprop_i),
        .l_TColl_2_1_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o),
        .l_TColl_2_1_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o_ap_vld),
        .l_TColl_0_2_0_constprop_i(l_TColl_0_2_0_constprop_i),
        .l_TColl_0_2_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o),
        .l_TColl_0_2_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o_ap_vld),
        .l_TColl_0_2_1_constprop_i(l_TColl_0_2_1_constprop_i),
        .l_TColl_0_2_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o),
        .l_TColl_0_2_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o_ap_vld),
        .l_TColl_0_2_2_constprop_i(l_TColl_0_2_2_constprop_i),
        .l_TColl_0_2_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o),
        .l_TColl_0_2_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o_ap_vld),
        .l_TColl_0_2_3_constprop_i(l_TColl_0_2_3_constprop_i),
        .l_TColl_0_2_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o),
        .l_TColl_0_2_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o_ap_vld),
        .l_TColl_1_2_0_constprop_i(l_TColl_1_2_0_constprop_i),
        .l_TColl_1_2_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o),
        .l_TColl_1_2_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o_ap_vld),
        .l_TColl_1_2_1_constprop_i(l_TColl_1_2_1_constprop_i),
        .l_TColl_1_2_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o),
        .l_TColl_1_2_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o_ap_vld),
        .l_TColl_1_2_2_constprop_i(l_TColl_1_2_2_constprop_i),
        .l_TColl_1_2_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o),
        .l_TColl_1_2_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o_ap_vld),
        .l_TColl_1_2_3_constprop_i(l_TColl_1_2_3_constprop_i),
        .l_TColl_1_2_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o),
        .l_TColl_1_2_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o_ap_vld),
        .l_TColl_2_2_0_constprop_i(l_TColl_2_2_0_constprop_i),
        .l_TColl_2_2_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o),
        .l_TColl_2_2_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o_ap_vld),
        .l_TColl_2_2_1_constprop_i(l_TColl_2_2_1_constprop_i),
        .l_TColl_2_2_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o),
        .l_TColl_2_2_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o_ap_vld),
        .l_TColl_2_2_2_constprop_i(l_TColl_2_2_2_constprop_i),
        .l_TColl_2_2_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o),
        .l_TColl_2_2_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o_ap_vld),
        .l_TColl_2_2_3_constprop_i(l_TColl_2_2_3_constprop_i),
        .l_TColl_2_2_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o),
        .l_TColl_2_2_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o_ap_vld),
        .l_TColl_0_3_0_constprop_i(l_TColl_0_3_0_constprop_i),
        .l_TColl_0_3_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o),
        .l_TColl_0_3_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o_ap_vld),
        .l_TColl_0_3_1_constprop_i(l_TColl_0_3_1_constprop_i),
        .l_TColl_0_3_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o),
        .l_TColl_0_3_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o_ap_vld),
        .l_TColl_0_3_2_constprop_i(l_TColl_0_3_2_constprop_i),
        .l_TColl_0_3_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o),
        .l_TColl_0_3_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o_ap_vld),
        .l_TColl_0_3_3_constprop_i(l_TColl_0_3_3_constprop_i),
        .l_TColl_0_3_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o),
        .l_TColl_0_3_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o_ap_vld),
        .l_TColl_1_3_0_constprop_i(l_TColl_1_3_0_constprop_i),
        .l_TColl_1_3_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o),
        .l_TColl_1_3_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o_ap_vld),
        .l_TColl_1_3_1_constprop_i(l_TColl_1_3_1_constprop_i),
        .l_TColl_1_3_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o),
        .l_TColl_1_3_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o_ap_vld),
        .l_TColl_1_3_2_constprop_i(l_TColl_1_3_2_constprop_i),
        .l_TColl_1_3_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o),
        .l_TColl_1_3_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o_ap_vld),
        .l_TColl_1_3_3_constprop_i(l_TColl_1_3_3_constprop_i),
        .l_TColl_1_3_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o),
        .l_TColl_1_3_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o_ap_vld),
        .l_TColl_2_3_0_constprop_i(l_TColl_2_3_0_constprop_i),
        .l_TColl_2_3_0_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o),
        .l_TColl_2_3_0_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o_ap_vld),
        .l_TColl_2_3_1_constprop_i(l_TColl_2_3_1_constprop_i),
        .l_TColl_2_3_1_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o),
        .l_TColl_2_3_1_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o_ap_vld),
        .l_TColl_2_3_2_constprop_i(l_TColl_2_3_2_constprop_i),
        .l_TColl_2_3_2_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o),
        .l_TColl_2_3_2_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o_ap_vld),
        .l_TColl_2_3_3_constprop_i(l_TColl_2_3_3_constprop_i),
        .l_TColl_2_3_3_constprop_o(grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o),
        .l_TColl_2_3_3_constprop_o_ap_vld(grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o_ap_vld),
        .ap_return(grp_detectCollNode_fu_1055_ap_return),
        .grp_fu_2529_p_din0(grp_detectCollNode_fu_1055_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_detectCollNode_fu_1055_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_detectCollNode_fu_1055_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_detectCollNode_fu_1055_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_detectCollNode_fu_1055_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_detectCollNode_fu_1055_grp_fu_2533_p_ce),
        .grp_fu_2537_p_din0(grp_detectCollNode_fu_1055_grp_fu_2537_p_din0),
        .grp_fu_2537_p_din1(grp_detectCollNode_fu_1055_grp_fu_2537_p_din1),
        .grp_fu_2537_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2537_p_opcode),
        .grp_fu_2537_p_dout0(grp_fu_2407_p_dout0),
        .grp_fu_2537_p_ce(grp_detectCollNode_fu_1055_grp_fu_2537_p_ce),
        .grp_fu_2541_p_din0(grp_detectCollNode_fu_1055_grp_fu_2541_p_din0),
        .grp_fu_2541_p_din1(grp_detectCollNode_fu_1055_grp_fu_2541_p_din1),
        .grp_fu_2541_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2541_p_opcode),
        .grp_fu_2541_p_dout0(grp_fu_2411_p_dout0),
        .grp_fu_2541_p_ce(grp_detectCollNode_fu_1055_grp_fu_2541_p_ce),
        .grp_fu_2545_p_din0(grp_detectCollNode_fu_1055_grp_fu_2545_p_din0),
        .grp_fu_2545_p_din1(grp_detectCollNode_fu_1055_grp_fu_2545_p_din1),
        .grp_fu_2545_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2545_p_opcode),
        .grp_fu_2545_p_dout0(grp_fu_2415_p_dout0),
        .grp_fu_2545_p_ce(grp_detectCollNode_fu_1055_grp_fu_2545_p_ce),
        .grp_fu_2549_p_din0(grp_detectCollNode_fu_1055_grp_fu_2549_p_din0),
        .grp_fu_2549_p_din1(grp_detectCollNode_fu_1055_grp_fu_2549_p_din1),
        .grp_fu_2549_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2549_p_opcode),
        .grp_fu_2549_p_dout0(grp_fu_2419_p_dout0),
        .grp_fu_2549_p_ce(grp_detectCollNode_fu_1055_grp_fu_2549_p_ce),
        .grp_fu_2553_p_din0(grp_detectCollNode_fu_1055_grp_fu_2553_p_din0),
        .grp_fu_2553_p_din1(grp_detectCollNode_fu_1055_grp_fu_2553_p_din1),
        .grp_fu_2553_p_opcode(grp_detectCollNode_fu_1055_grp_fu_2553_p_opcode),
        .grp_fu_2553_p_dout0(grp_fu_2423_p_dout0),
        .grp_fu_2553_p_ce(grp_detectCollNode_fu_1055_grp_fu_2553_p_ce),
        .grp_fu_2557_p_din0(grp_detectCollNode_fu_1055_grp_fu_2557_p_din0),
        .grp_fu_2557_p_din1(grp_detectCollNode_fu_1055_grp_fu_2557_p_din1),
        .grp_fu_2557_p_dout0(grp_fu_2435_p_dout0),
        .grp_fu_2557_p_ce(grp_detectCollNode_fu_1055_grp_fu_2557_p_ce),
        .grp_fu_2561_p_din0(grp_detectCollNode_fu_1055_grp_fu_2561_p_din0),
        .grp_fu_2561_p_din1(grp_detectCollNode_fu_1055_grp_fu_2561_p_din1),
        .grp_fu_2561_p_dout0(grp_fu_2439_p_dout0),
        .grp_fu_2561_p_ce(grp_detectCollNode_fu_1055_grp_fu_2561_p_ce),
        .grp_fu_2565_p_din0(grp_detectCollNode_fu_1055_grp_fu_2565_p_din0),
        .grp_fu_2565_p_din1(grp_detectCollNode_fu_1055_grp_fu_2565_p_din1),
        .grp_fu_2565_p_dout0(grp_fu_2443_p_dout0),
        .grp_fu_2565_p_ce(grp_detectCollNode_fu_1055_grp_fu_2565_p_ce),
        .grp_fu_1454_p_din0(grp_detectCollNode_fu_1055_grp_fu_1454_p_din0),
        .grp_fu_1454_p_din1(grp_detectCollNode_fu_1055_grp_fu_1454_p_din1),
        .grp_fu_1454_p_opcode(grp_detectCollNode_fu_1055_grp_fu_1454_p_opcode),
        .grp_fu_1454_p_dout0(grp_fu_1454_p2),
        .grp_fu_1454_p_ce(grp_detectCollNode_fu_1055_grp_fu_1454_p_ce),
        .grp_fu_1462_p_din0(grp_detectCollNode_fu_1055_grp_fu_1462_p_din0),
        .grp_fu_1462_p_din1(grp_detectCollNode_fu_1055_grp_fu_1462_p_din1),
        .grp_fu_1462_p_dout0(grp_fu_1462_p2),
        .grp_fu_1462_p_ce(grp_detectCollNode_fu_1055_grp_fu_1462_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_293_19 grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_ready),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .dist_6_out(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_dist_6_out),
        .dist_6_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_dist_6_out_ap_vld),
        .goal_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_address0),
        .goal_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_ce0),
        .goal_q0(goal_q0),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110 grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404(
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_ready),
        .minDist_4(reg_1470),
        .sub_ln296_1(sub_ln296_1_reg_2498),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .bestIdx_6_out(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out),
        .bestIdx_6_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out_ap_vld),
        .goal_address0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_address0),
        .goal_ce0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_ce0),
        .goal_q0(goal_q0),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_ce),
        .grp_fu_1454_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din0),
        .grp_fu_1454_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din1),
        .grp_fu_1454_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_opcode),
        .grp_fu_1454_p_dout0(grp_fu_1454_p2),
        .grp_fu_1454_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_ce),
        .grp_fu_1462_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din0),
        .grp_fu_1462_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din1),
        .grp_fu_1462_p_dout0(grp_fu_1462_p2),
        .grp_fu_1462_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_293_111 grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_ready),
        .sub_ln294_1(sub_ln294_reg_2503),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_ce0),
        .rrtVertices_q0(rrtVertices_q0),
        .dist_10_out(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_dist_10_out),
        .dist_10_out_ap_vld(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_dist_10_out_ap_vld),
        .goal_address0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_address0),
        .goal_ce0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_ce0),
        .goal_q0(goal_q0),
        .grp_fu_2529_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din0),
        .grp_fu_2529_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din1),
        .grp_fu_2529_p_opcode(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_opcode),
        .grp_fu_2529_p_dout0(grp_fu_2403_p_dout0),
        .grp_fu_2529_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_ce),
        .grp_fu_2533_p_din0(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din0),
        .grp_fu_2533_p_din1(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din1),
        .grp_fu_2533_p_dout0(grp_fu_2431_p_dout0),
        .grp_fu_2533_p_ce(grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_ce)
    );

    main_planRRT_Pipeline_VITIS_LOOP_139_9 grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start),
        .ap_done(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_done),
        .ap_idle(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_idle),
        .ap_ready(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_ready),
        .sub_ln139(sub_ln139_reg_2524),
        .rrtVertices_address0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_address0),
        .rrtVertices_ce0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_ce0),
        .rrtVertices_we0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_we0),
        .rrtVertices_d0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_d0),
        .goal_address0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_address0),
        .goal_ce0(grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_ce0),
        .goal_q0(goal_q0)
    );

    main_fmul_32ns_32ns_32_4_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fmul_32ns_32ns_32_4_max_dsp_1_U1611 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1431_p0),
        .din1(grp_fu_1431_p1),
        .ce(grp_fu_1431_ce),
        .dout(grp_fu_1431_p2)
    );

    main_uitofp_32ns_32_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(32)
    ) uitofp_32ns_32_6_no_dsp_1_U1612 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1436_p0),
        .ce(grp_fu_1436_ce),
        .dout(grp_fu_1436_p1)
    );

    main_fpext_32ns_64_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) fpext_32ns_64_2_no_dsp_1_U1613 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1439_p0),
        .ce(grp_fu_1439_ce),
        .dout(grp_fu_1439_p1)
    );

    main_ddiv_64ns_64ns_64_59_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(59),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) ddiv_64ns_64ns_64_59_no_dsp_1_U1615 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(64'd4598175219545276416),
        .din1(reg_1470),
        .ce(1'b1),
        .dout(grp_fu_1448_p2)
    );

    main_dcmp_64ns_64ns_1_2_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(1)
    ) dcmp_64ns_64ns_1_2_no_dsp_1_U1616 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1454_p0),
        .din1(grp_fu_1454_p1),
        .ce(grp_fu_1454_ce),
        .opcode(grp_fu_1454_opcode),
        .dout(grp_fu_1454_p2)
    );

    main_dsqrt_64ns_64ns_64_57_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(57),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dsqrt_64ns_64ns_64_57_no_dsp_1_U1617 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_1462_p0),
        .din1(grp_fu_1462_p1),
        .ce(grp_fu_1462_ce),
        .dout(grp_fu_1462_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_detectCollNode_fu_1055_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state208)) begin
                grp_detectCollNode_fu_1055_ap_start_reg <= 1'b1;
            end else if ((grp_detectCollNode_fu_1055_ap_ready == 1'b1)) begin
                grp_detectCollNode_fu_1055_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd1 == and_ln110_fu_1614_p2) & (1'b1 == ap_CS_fsm_state19))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state82)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state203)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd0 == and_ln119_fu_1767_p2) & (1'b1 == ap_CS_fsm_state144))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd0 == and_ln188_fu_1809_p2) & (1'b1 == ap_CS_fsm_state206))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd1 == and_ln138_fu_1960_p2) & (1'b1 == ap_CS_fsm_state337))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state3) & (icmp_ln107_fu_1491_p2 == 1'd1))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg <= 1'b0;
        end else begin
            if (((1'd1 == and_ln188_fu_1809_p2) & (1'b1 == ap_CS_fsm_state206))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state277)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state84)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_state209_on_subcall_done) & (1'b1 == ap_CS_fsm_state209) & ((1'd0 == and_ln188_reg_2467) | (grp_detectCollNode_fu_1055_ap_return == 1'd1)))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state21)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg <= 1'b0;
        end else begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state275)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state80)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg <= 1'b1;
            end else if ((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_ready == 1'b1)) begin
                grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            numVertices_fu_520 <= 32'd1;
        end else if (((1'b1 == ap_CS_fsm_state216) & (grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_done == 1'b1))) begin
            numVertices_fu_520 <= numVertices_2_fu_1815_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state215)) begin
            s_reg_960 <= grp_fu_2427_p_dout0;
        end else if (((1'b0 == ap_block_state204_on_subcall_done) & (1'b1 == ap_CS_fsm_state204))) begin
            s_reg_960 <= 64'd0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state19)) begin
            and_ln110_reg_2427 <= and_ln110_fu_1614_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state144)) begin
            and_ln119_reg_2458 <= and_ln119_fu_1767_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state206)) begin
            and_ln188_reg_2467 <= and_ln188_fu_1809_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state81) & (grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out_ap_vld == 1'b1))) begin
            bestIdx_3_loc_fu_540 <= grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_bestIdx_3_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state276))) begin
            bestIdx_6_loc_fu_528 <= grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_bestIdx_6_out;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state11)) begin
            conv_i1_reg_2401 <= grp_fu_1436_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state17)) begin
            conv_reg_2411 <= grp_fu_1439_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state15)) begin
            div_i_reg_2406 <= grp_fu_1431_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state203)) begin
            f_reg_2462 <= grp_fu_1448_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            icmp_ln107_reg_2379 <= icmp_ln107_fu_1491_p2;
            numVertices_1_reg_2362 <= numVertices_fu_520;
            trunc_ln83_1_reg_2374 <= trunc_ln83_1_fu_1487_p1;
            trunc_ln83_reg_2369 <= trunc_ln83_fu_1483_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state18)) begin
            icmp_ln110_1_reg_2422 <= icmp_ln110_1_fu_1604_p2;
            icmp_ln110_reg_2417   <= icmp_ln110_fu_1598_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state336)) begin
            icmp_ln138_1_reg_2516 <= icmp_ln138_1_fu_1950_p2;
            icmp_ln138_reg_2511   <= icmp_ln138_fu_1944_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state6)) begin
            lfsr <= rand_int_fu_1564_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            lshr_ln_reg_2386 <= {
                {grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out[15:1]}
            };
            xor_ln38_reg_2391 <= xor_ln38_fu_1558_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state335) | (1'b1 == ap_CS_fsm_state274) | (1'b1 == ap_CS_fsm_state142) | (1'b1 == ap_CS_fsm_state79))) begin
            reg_1470 <= grp_fu_1462_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state274)) begin
            select_ln96_5_reg_2492 <= select_ln96_5_fu_1859_p3;
            trunc_ln83_2_reg_2482  <= trunc_ln83_2_fu_1829_p1;
            trunc_ln83_3_reg_2487  <= trunc_ln83_3_fu_1833_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state79)) begin
            select_ln96_reg_2439 <= select_ln96_fu_1664_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state82)) begin
            sub_ln114_reg_2450[12 : 1] <= sub_ln114_fu_1720_p2[12 : 1];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state20)) begin
            sub_ln130_reg_2431[12 : 1] <= sub_ln130_fu_1634_p2[12 : 1];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state337)) begin
            sub_ln139_reg_2524[12 : 1] <= sub_ln139_fu_1980_p2[12 : 1];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state277)) begin
            sub_ln294_reg_2503[12 : 1] <= sub_ln294_fu_1915_p2[12 : 1];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state275)) begin
            sub_ln296_1_reg_2498[34 : 1] <= sub_ln296_1_fu_1885_p2[34 : 1];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state80)) begin
            sub_ln296_reg_2445[34 : 1] <= sub_ln296_fu_1690_p2[34 : 1];
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (1'b1 == ap_CS_fsm_state209))) begin
            ang_address0 = grp_detectCollNode_fu_1055_ang_address0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            ang_address0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_address0;
        end else begin
            ang_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (1'b1 == ap_CS_fsm_state209))) begin
            ang_ce0 = grp_detectCollNode_fu_1055_ang_ce0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            ang_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_ce0;
        end else begin
            ang_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state207)) begin
            ang_we0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ang_we0;
        end else begin
            ang_we0 = 1'b0;
        end
    end

    assign ap_ST_fsm_state100_blk = 1'b0;

    assign ap_ST_fsm_state101_blk = 1'b0;

    assign ap_ST_fsm_state102_blk = 1'b0;

    assign ap_ST_fsm_state103_blk = 1'b0;

    assign ap_ST_fsm_state104_blk = 1'b0;

    assign ap_ST_fsm_state105_blk = 1'b0;

    assign ap_ST_fsm_state106_blk = 1'b0;

    assign ap_ST_fsm_state107_blk = 1'b0;

    assign ap_ST_fsm_state108_blk = 1'b0;

    assign ap_ST_fsm_state109_blk = 1'b0;

    assign ap_ST_fsm_state10_blk  = 1'b0;

    assign ap_ST_fsm_state110_blk = 1'b0;

    assign ap_ST_fsm_state111_blk = 1'b0;

    assign ap_ST_fsm_state112_blk = 1'b0;

    assign ap_ST_fsm_state113_blk = 1'b0;

    assign ap_ST_fsm_state114_blk = 1'b0;

    assign ap_ST_fsm_state115_blk = 1'b0;

    assign ap_ST_fsm_state116_blk = 1'b0;

    assign ap_ST_fsm_state117_blk = 1'b0;

    assign ap_ST_fsm_state118_blk = 1'b0;

    assign ap_ST_fsm_state119_blk = 1'b0;

    assign ap_ST_fsm_state11_blk  = 1'b0;

    assign ap_ST_fsm_state120_blk = 1'b0;

    assign ap_ST_fsm_state121_blk = 1'b0;

    assign ap_ST_fsm_state122_blk = 1'b0;

    assign ap_ST_fsm_state123_blk = 1'b0;

    assign ap_ST_fsm_state124_blk = 1'b0;

    assign ap_ST_fsm_state125_blk = 1'b0;

    assign ap_ST_fsm_state126_blk = 1'b0;

    assign ap_ST_fsm_state127_blk = 1'b0;

    assign ap_ST_fsm_state128_blk = 1'b0;

    assign ap_ST_fsm_state129_blk = 1'b0;

    assign ap_ST_fsm_state12_blk  = 1'b0;

    assign ap_ST_fsm_state130_blk = 1'b0;

    assign ap_ST_fsm_state131_blk = 1'b0;

    assign ap_ST_fsm_state132_blk = 1'b0;

    assign ap_ST_fsm_state133_blk = 1'b0;

    assign ap_ST_fsm_state134_blk = 1'b0;

    assign ap_ST_fsm_state135_blk = 1'b0;

    assign ap_ST_fsm_state136_blk = 1'b0;

    assign ap_ST_fsm_state137_blk = 1'b0;

    assign ap_ST_fsm_state138_blk = 1'b0;

    assign ap_ST_fsm_state139_blk = 1'b0;

    assign ap_ST_fsm_state13_blk  = 1'b0;

    assign ap_ST_fsm_state140_blk = 1'b0;

    assign ap_ST_fsm_state141_blk = 1'b0;

    assign ap_ST_fsm_state142_blk = 1'b0;

    assign ap_ST_fsm_state143_blk = 1'b0;

    assign ap_ST_fsm_state144_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_done == 1'b0)) begin
            ap_ST_fsm_state145_blk = 1'b1;
        end else begin
            ap_ST_fsm_state145_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state146_blk = 1'b0;

    assign ap_ST_fsm_state147_blk = 1'b0;

    assign ap_ST_fsm_state148_blk = 1'b0;

    assign ap_ST_fsm_state149_blk = 1'b0;

    assign ap_ST_fsm_state14_blk  = 1'b0;

    assign ap_ST_fsm_state150_blk = 1'b0;

    assign ap_ST_fsm_state151_blk = 1'b0;

    assign ap_ST_fsm_state152_blk = 1'b0;

    assign ap_ST_fsm_state153_blk = 1'b0;

    assign ap_ST_fsm_state154_blk = 1'b0;

    assign ap_ST_fsm_state155_blk = 1'b0;

    assign ap_ST_fsm_state156_blk = 1'b0;

    assign ap_ST_fsm_state157_blk = 1'b0;

    assign ap_ST_fsm_state158_blk = 1'b0;

    assign ap_ST_fsm_state159_blk = 1'b0;

    assign ap_ST_fsm_state15_blk  = 1'b0;

    assign ap_ST_fsm_state160_blk = 1'b0;

    assign ap_ST_fsm_state161_blk = 1'b0;

    assign ap_ST_fsm_state162_blk = 1'b0;

    assign ap_ST_fsm_state163_blk = 1'b0;

    assign ap_ST_fsm_state164_blk = 1'b0;

    assign ap_ST_fsm_state165_blk = 1'b0;

    assign ap_ST_fsm_state166_blk = 1'b0;

    assign ap_ST_fsm_state167_blk = 1'b0;

    assign ap_ST_fsm_state168_blk = 1'b0;

    assign ap_ST_fsm_state169_blk = 1'b0;

    assign ap_ST_fsm_state16_blk  = 1'b0;

    assign ap_ST_fsm_state170_blk = 1'b0;

    assign ap_ST_fsm_state171_blk = 1'b0;

    assign ap_ST_fsm_state172_blk = 1'b0;

    assign ap_ST_fsm_state173_blk = 1'b0;

    assign ap_ST_fsm_state174_blk = 1'b0;

    assign ap_ST_fsm_state175_blk = 1'b0;

    assign ap_ST_fsm_state176_blk = 1'b0;

    assign ap_ST_fsm_state177_blk = 1'b0;

    assign ap_ST_fsm_state178_blk = 1'b0;

    assign ap_ST_fsm_state179_blk = 1'b0;

    assign ap_ST_fsm_state17_blk  = 1'b0;

    assign ap_ST_fsm_state180_blk = 1'b0;

    assign ap_ST_fsm_state181_blk = 1'b0;

    assign ap_ST_fsm_state182_blk = 1'b0;

    assign ap_ST_fsm_state183_blk = 1'b0;

    assign ap_ST_fsm_state184_blk = 1'b0;

    assign ap_ST_fsm_state185_blk = 1'b0;

    assign ap_ST_fsm_state186_blk = 1'b0;

    assign ap_ST_fsm_state187_blk = 1'b0;

    assign ap_ST_fsm_state188_blk = 1'b0;

    assign ap_ST_fsm_state189_blk = 1'b0;

    assign ap_ST_fsm_state18_blk  = 1'b0;

    assign ap_ST_fsm_state190_blk = 1'b0;

    assign ap_ST_fsm_state191_blk = 1'b0;

    assign ap_ST_fsm_state192_blk = 1'b0;

    assign ap_ST_fsm_state193_blk = 1'b0;

    assign ap_ST_fsm_state194_blk = 1'b0;

    assign ap_ST_fsm_state195_blk = 1'b0;

    assign ap_ST_fsm_state196_blk = 1'b0;

    assign ap_ST_fsm_state197_blk = 1'b0;

    assign ap_ST_fsm_state198_blk = 1'b0;

    assign ap_ST_fsm_state199_blk = 1'b0;

    assign ap_ST_fsm_state19_blk  = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state200_blk = 1'b0;

    assign ap_ST_fsm_state201_blk = 1'b0;

    assign ap_ST_fsm_state202_blk = 1'b0;

    assign ap_ST_fsm_state203_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state204_on_subcall_done)) begin
            ap_ST_fsm_state204_blk = 1'b1;
        end else begin
            ap_ST_fsm_state204_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state205_blk = 1'b0;

    assign ap_ST_fsm_state206_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_done == 1'b0)) begin
            ap_ST_fsm_state207_blk = 1'b1;
        end else begin
            ap_ST_fsm_state207_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state208_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state209_on_subcall_done)) begin
            ap_ST_fsm_state209_blk = 1'b1;
        end else begin
            ap_ST_fsm_state209_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_block_state20_on_subcall_done)) begin
            ap_ST_fsm_state20_blk = 1'b1;
        end else begin
            ap_ST_fsm_state20_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state210_blk = 1'b0;

    assign ap_ST_fsm_state211_blk = 1'b0;

    assign ap_ST_fsm_state212_blk = 1'b0;

    assign ap_ST_fsm_state213_blk = 1'b0;

    assign ap_ST_fsm_state214_blk = 1'b0;

    assign ap_ST_fsm_state215_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_done == 1'b0)) begin
            ap_ST_fsm_state216_blk = 1'b1;
        end else begin
            ap_ST_fsm_state216_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_done == 1'b0)) begin
            ap_ST_fsm_state217_blk = 1'b1;
        end else begin
            ap_ST_fsm_state217_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state218_blk = 1'b0;

    assign ap_ST_fsm_state219_blk = 1'b0;

    assign ap_ST_fsm_state21_blk  = 1'b0;

    assign ap_ST_fsm_state220_blk = 1'b0;

    assign ap_ST_fsm_state221_blk = 1'b0;

    assign ap_ST_fsm_state222_blk = 1'b0;

    assign ap_ST_fsm_state223_blk = 1'b0;

    assign ap_ST_fsm_state224_blk = 1'b0;

    assign ap_ST_fsm_state225_blk = 1'b0;

    assign ap_ST_fsm_state226_blk = 1'b0;

    assign ap_ST_fsm_state227_blk = 1'b0;

    assign ap_ST_fsm_state228_blk = 1'b0;

    assign ap_ST_fsm_state229_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_done == 1'b0)) begin
            ap_ST_fsm_state22_blk = 1'b1;
        end else begin
            ap_ST_fsm_state22_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state230_blk = 1'b0;

    assign ap_ST_fsm_state231_blk = 1'b0;

    assign ap_ST_fsm_state232_blk = 1'b0;

    assign ap_ST_fsm_state233_blk = 1'b0;

    assign ap_ST_fsm_state234_blk = 1'b0;

    assign ap_ST_fsm_state235_blk = 1'b0;

    assign ap_ST_fsm_state236_blk = 1'b0;

    assign ap_ST_fsm_state237_blk = 1'b0;

    assign ap_ST_fsm_state238_blk = 1'b0;

    assign ap_ST_fsm_state239_blk = 1'b0;

    assign ap_ST_fsm_state23_blk  = 1'b0;

    assign ap_ST_fsm_state240_blk = 1'b0;

    assign ap_ST_fsm_state241_blk = 1'b0;

    assign ap_ST_fsm_state242_blk = 1'b0;

    assign ap_ST_fsm_state243_blk = 1'b0;

    assign ap_ST_fsm_state244_blk = 1'b0;

    assign ap_ST_fsm_state245_blk = 1'b0;

    assign ap_ST_fsm_state246_blk = 1'b0;

    assign ap_ST_fsm_state247_blk = 1'b0;

    assign ap_ST_fsm_state248_blk = 1'b0;

    assign ap_ST_fsm_state249_blk = 1'b0;

    assign ap_ST_fsm_state24_blk  = 1'b0;

    assign ap_ST_fsm_state250_blk = 1'b0;

    assign ap_ST_fsm_state251_blk = 1'b0;

    assign ap_ST_fsm_state252_blk = 1'b0;

    assign ap_ST_fsm_state253_blk = 1'b0;

    assign ap_ST_fsm_state254_blk = 1'b0;

    assign ap_ST_fsm_state255_blk = 1'b0;

    assign ap_ST_fsm_state256_blk = 1'b0;

    assign ap_ST_fsm_state257_blk = 1'b0;

    assign ap_ST_fsm_state258_blk = 1'b0;

    assign ap_ST_fsm_state259_blk = 1'b0;

    assign ap_ST_fsm_state25_blk  = 1'b0;

    assign ap_ST_fsm_state260_blk = 1'b0;

    assign ap_ST_fsm_state261_blk = 1'b0;

    assign ap_ST_fsm_state262_blk = 1'b0;

    assign ap_ST_fsm_state263_blk = 1'b0;

    assign ap_ST_fsm_state264_blk = 1'b0;

    assign ap_ST_fsm_state265_blk = 1'b0;

    assign ap_ST_fsm_state266_blk = 1'b0;

    assign ap_ST_fsm_state267_blk = 1'b0;

    assign ap_ST_fsm_state268_blk = 1'b0;

    assign ap_ST_fsm_state269_blk = 1'b0;

    assign ap_ST_fsm_state26_blk  = 1'b0;

    assign ap_ST_fsm_state270_blk = 1'b0;

    assign ap_ST_fsm_state271_blk = 1'b0;

    assign ap_ST_fsm_state272_blk = 1'b0;

    assign ap_ST_fsm_state273_blk = 1'b0;

    assign ap_ST_fsm_state274_blk = 1'b0;

    assign ap_ST_fsm_state275_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_done == 1'b0)) begin
            ap_ST_fsm_state276_blk = 1'b1;
        end else begin
            ap_ST_fsm_state276_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state277_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_done == 1'b0)) begin
            ap_ST_fsm_state278_blk = 1'b1;
        end else begin
            ap_ST_fsm_state278_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state279_blk = 1'b0;

    assign ap_ST_fsm_state27_blk  = 1'b0;

    assign ap_ST_fsm_state280_blk = 1'b0;

    assign ap_ST_fsm_state281_blk = 1'b0;

    assign ap_ST_fsm_state282_blk = 1'b0;

    assign ap_ST_fsm_state283_blk = 1'b0;

    assign ap_ST_fsm_state284_blk = 1'b0;

    assign ap_ST_fsm_state285_blk = 1'b0;

    assign ap_ST_fsm_state286_blk = 1'b0;

    assign ap_ST_fsm_state287_blk = 1'b0;

    assign ap_ST_fsm_state288_blk = 1'b0;

    assign ap_ST_fsm_state289_blk = 1'b0;

    assign ap_ST_fsm_state28_blk  = 1'b0;

    assign ap_ST_fsm_state290_blk = 1'b0;

    assign ap_ST_fsm_state291_blk = 1'b0;

    assign ap_ST_fsm_state292_blk = 1'b0;

    assign ap_ST_fsm_state293_blk = 1'b0;

    assign ap_ST_fsm_state294_blk = 1'b0;

    assign ap_ST_fsm_state295_blk = 1'b0;

    assign ap_ST_fsm_state296_blk = 1'b0;

    assign ap_ST_fsm_state297_blk = 1'b0;

    assign ap_ST_fsm_state298_blk = 1'b0;

    assign ap_ST_fsm_state299_blk = 1'b0;

    assign ap_ST_fsm_state29_blk  = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_done == 1'b0)) begin
            ap_ST_fsm_state2_blk = 1'b1;
        end else begin
            ap_ST_fsm_state2_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state300_blk = 1'b0;

    assign ap_ST_fsm_state301_blk = 1'b0;

    assign ap_ST_fsm_state302_blk = 1'b0;

    assign ap_ST_fsm_state303_blk = 1'b0;

    assign ap_ST_fsm_state304_blk = 1'b0;

    assign ap_ST_fsm_state305_blk = 1'b0;

    assign ap_ST_fsm_state306_blk = 1'b0;

    assign ap_ST_fsm_state307_blk = 1'b0;

    assign ap_ST_fsm_state308_blk = 1'b0;

    assign ap_ST_fsm_state309_blk = 1'b0;

    assign ap_ST_fsm_state30_blk  = 1'b0;

    assign ap_ST_fsm_state310_blk = 1'b0;

    assign ap_ST_fsm_state311_blk = 1'b0;

    assign ap_ST_fsm_state312_blk = 1'b0;

    assign ap_ST_fsm_state313_blk = 1'b0;

    assign ap_ST_fsm_state314_blk = 1'b0;

    assign ap_ST_fsm_state315_blk = 1'b0;

    assign ap_ST_fsm_state316_blk = 1'b0;

    assign ap_ST_fsm_state317_blk = 1'b0;

    assign ap_ST_fsm_state318_blk = 1'b0;

    assign ap_ST_fsm_state319_blk = 1'b0;

    assign ap_ST_fsm_state31_blk  = 1'b0;

    assign ap_ST_fsm_state320_blk = 1'b0;

    assign ap_ST_fsm_state321_blk = 1'b0;

    assign ap_ST_fsm_state322_blk = 1'b0;

    assign ap_ST_fsm_state323_blk = 1'b0;

    assign ap_ST_fsm_state324_blk = 1'b0;

    assign ap_ST_fsm_state325_blk = 1'b0;

    assign ap_ST_fsm_state326_blk = 1'b0;

    assign ap_ST_fsm_state327_blk = 1'b0;

    assign ap_ST_fsm_state328_blk = 1'b0;

    assign ap_ST_fsm_state329_blk = 1'b0;

    assign ap_ST_fsm_state32_blk  = 1'b0;

    assign ap_ST_fsm_state330_blk = 1'b0;

    assign ap_ST_fsm_state331_blk = 1'b0;

    assign ap_ST_fsm_state332_blk = 1'b0;

    assign ap_ST_fsm_state333_blk = 1'b0;

    assign ap_ST_fsm_state334_blk = 1'b0;

    assign ap_ST_fsm_state335_blk = 1'b0;

    assign ap_ST_fsm_state336_blk = 1'b0;

    assign ap_ST_fsm_state337_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state338_on_subcall_done)) begin
            ap_ST_fsm_state338_blk = 1'b1;
        end else begin
            ap_ST_fsm_state338_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_done == 1'b0)) begin
            ap_ST_fsm_state4_blk = 1'b1;
        end else begin
            ap_ST_fsm_state4_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    assign ap_ST_fsm_state73_blk = 1'b0;

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state75_blk = 1'b0;

    assign ap_ST_fsm_state76_blk = 1'b0;

    assign ap_ST_fsm_state77_blk = 1'b0;

    assign ap_ST_fsm_state78_blk = 1'b0;

    assign ap_ST_fsm_state79_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state80_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_done == 1'b0)) begin
            ap_ST_fsm_state81_blk = 1'b1;
        end else begin
            ap_ST_fsm_state81_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state82_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_done == 1'b0)) begin
            ap_ST_fsm_state83_blk = 1'b1;
        end else begin
            ap_ST_fsm_state83_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state84_blk = 1'b0;

    always @(*) begin
        if ((grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_done == 1'b0)) begin
            ap_ST_fsm_state85_blk = 1'b1;
        end else begin
            ap_ST_fsm_state85_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state86_blk = 1'b0;

    assign ap_ST_fsm_state87_blk = 1'b0;

    assign ap_ST_fsm_state88_blk = 1'b0;

    assign ap_ST_fsm_state89_blk = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state90_blk = 1'b0;

    assign ap_ST_fsm_state91_blk = 1'b0;

    assign ap_ST_fsm_state92_blk = 1'b0;

    assign ap_ST_fsm_state93_blk = 1'b0;

    assign ap_ST_fsm_state94_blk = 1'b0;

    assign ap_ST_fsm_state95_blk = 1'b0;

    assign ap_ST_fsm_state96_blk = 1'b0;

    assign ap_ST_fsm_state97_blk = 1'b0;

    assign ap_ST_fsm_state98_blk = 1'b0;

    assign ap_ST_fsm_state99_blk = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if ((((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) | ((1'b0 == ap_block_state338_on_subcall_done) & (1'b1 == ap_CS_fsm_state338)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_state338_on_subcall_done) & (1'b1 == ap_CS_fsm_state338))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            goal_address0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_address0;
        end else if ((1'b1 == ap_CS_fsm_state278)) begin
            goal_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_address0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            goal_address0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_address0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            goal_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_address0;
        end else if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            goal_address0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_address0;
        end else begin
            goal_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            goal_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_goal_ce0;
        end else if ((1'b1 == ap_CS_fsm_state278)) begin
            goal_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_goal_ce0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            goal_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_goal_ce0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            goal_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_goal_ce0;
        end else if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            goal_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_goal_ce0;
        end else begin
            goal_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1431_ce = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_ce;
        end else begin
            grp_fu_1431_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1431_p0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_1431_p0 = conv_i1_reg_2401;
        end else begin
            grp_fu_1431_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1431_p1 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1431_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_fu_1431_p1 = 32'd796917760;
        end else begin
            grp_fu_1431_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1436_ce = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_ce;
        end else begin
            grp_fu_1436_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1436_p0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1436_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            grp_fu_1436_p0 = zext_ln47_fu_1576_p1;
        end else begin
            grp_fu_1436_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1439_ce = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_ce;
        end else begin
            grp_fu_1439_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_1439_p0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_1439_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state16)) begin
            grp_fu_1439_p0 = div_i_reg_2406;
        end else begin
            grp_fu_1439_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state214) | (1'b1 == ap_CS_fsm_state213) | (1'b1 == ap_CS_fsm_state212) | (1'b1 == ap_CS_fsm_state211) | (1'b1 == ap_CS_fsm_state210) | (1'b1 == ap_CS_fsm_state215) | ((1'b0 == ap_block_state209_on_subcall_done) & (1'b1 == ap_CS_fsm_state209)))) begin
            grp_fu_1442_ce = 1'b1;
        end else begin
            grp_fu_1442_ce = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1454_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1454_ce = grp_detectCollNode_fu_1055_grp_fu_1454_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1454_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_ce;
        end else begin
            grp_fu_1454_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1454_opcode = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1454_opcode = grp_detectCollNode_fu_1055_grp_fu_1454_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1454_opcode = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state205)) begin
            grp_fu_1454_opcode = 5'd5;
        end else if ((1'b1 == ap_CS_fsm_state143)) begin
            grp_fu_1454_opcode = 5'd2;
        end else if (((1'b1 == ap_CS_fsm_state336) | (1'b1 == ap_CS_fsm_state18))) begin
            grp_fu_1454_opcode = 5'd4;
        end else begin
            grp_fu_1454_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1454_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1454_p0 = grp_detectCollNode_fu_1055_grp_fu_1454_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1454_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state205)) begin
            grp_fu_1454_p0 = s_reg_960;
        end else if (((1'b1 == ap_CS_fsm_state143) | (1'b1 == ap_CS_fsm_state336))) begin
            grp_fu_1454_p0 = reg_1470;
        end else if ((1'b1 == ap_CS_fsm_state18)) begin
            grp_fu_1454_p0 = conv_reg_2411;
        end else begin
            grp_fu_1454_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1454_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1454_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1454_p1 = grp_detectCollNode_fu_1055_grp_fu_1454_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1454_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1454_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state205)) begin
            grp_fu_1454_p1 = 64'd4607182418800017408;
        end else if (((1'b1 == ap_CS_fsm_state143) | (1'b1 == ap_CS_fsm_state336))) begin
            grp_fu_1454_p1 = 64'd4598175219545276416;
        end else if ((1'b1 == ap_CS_fsm_state18)) begin
            grp_fu_1454_p1 = 64'd4587366580439587226;
        end else begin
            grp_fu_1454_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1462_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1462_ce = grp_detectCollNode_fu_1055_grp_fu_1462_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1462_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_ce;
        end else begin
            grp_fu_1462_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1462_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1462_p0 = grp_detectCollNode_fu_1055_grp_fu_1462_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1462_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din0;
        end else begin
            grp_fu_1462_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_1462_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_1462_p1 = grp_detectCollNode_fu_1055_grp_fu_1462_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_1462_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state279)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_dist_10_out;
        end else if ((1'b1 == ap_CS_fsm_state218)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_dist_6_out;
        end else if ((1'b1 == ap_CS_fsm_state86)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_dist_4_out;
        end else if ((1'b1 == ap_CS_fsm_state23)) begin
            grp_fu_1462_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_dist_out;
        end else begin
            grp_fu_1462_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2529_ce = grp_detectCollNode_fu_1055_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2529_ce = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_ce;
        end else begin
            grp_fu_2529_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2529_opcode = grp_detectCollNode_fu_1055_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2529_opcode = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_opcode;
        end else begin
            grp_fu_2529_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2529_p0 = grp_detectCollNode_fu_1055_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2529_p0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din0;
        end else begin
            grp_fu_2529_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2529_p1 = grp_detectCollNode_fu_1055_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2529_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2529_p1 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2529_p_din1;
        end else begin
            grp_fu_2529_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2533_ce = grp_detectCollNode_fu_1055_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2533_ce = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_ce;
        end else begin
            grp_fu_2533_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2533_p0 = grp_detectCollNode_fu_1055_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2533_p0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din0;
        end else begin
            grp_fu_2533_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state278)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2533_p1 = grp_detectCollNode_fu_1055_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_grp_fu_2533_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_2533_p1 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_grp_fu_2533_p_din1;
        end else begin
            grp_fu_2533_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2537_ce = grp_detectCollNode_fu_1055_grp_fu_2537_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2537_ce = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_ce;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2537_ce = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_ce;
        end else begin
            grp_fu_2537_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2537_opcode = grp_detectCollNode_fu_1055_grp_fu_2537_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2537_opcode = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_opcode;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2537_opcode = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_opcode;
        end else begin
            grp_fu_2537_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2537_p0 = grp_detectCollNode_fu_1055_grp_fu_2537_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2537_p0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din0;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2537_p0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din0;
        end else begin
            grp_fu_2537_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2537_p1 = grp_detectCollNode_fu_1055_grp_fu_2537_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            grp_fu_2537_p1 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_grp_fu_2537_p_din1;
        end else if ((1'b1 == ap_CS_fsm_state204)) begin
            grp_fu_2537_p1 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_grp_fu_2537_p_din1;
        end else begin
            grp_fu_2537_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2541_ce = grp_detectCollNode_fu_1055_grp_fu_2541_p_ce;
        end else begin
            grp_fu_2541_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2545_ce = grp_detectCollNode_fu_1055_grp_fu_2545_p_ce;
        end else begin
            grp_fu_2545_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2549_ce = grp_detectCollNode_fu_1055_grp_fu_2549_p_ce;
        end else begin
            grp_fu_2549_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2553_ce = grp_detectCollNode_fu_1055_grp_fu_2553_p_ce;
        end else begin
            grp_fu_2553_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2557_ce = grp_detectCollNode_fu_1055_grp_fu_2557_p_ce;
        end else begin
            grp_fu_2557_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2561_ce = grp_detectCollNode_fu_1055_grp_fu_2561_p_ce;
        end else begin
            grp_fu_2561_ce = 1'b1;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state209)) begin
            grp_fu_2565_ce = grp_detectCollNode_fu_1055_grp_fu_2565_p_ce;
        end else begin
            grp_fu_2565_ce = 1'b1;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_0_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o;
        end else begin
            l_TColl_0_0_0_constprop_o = l_TColl_0_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_0_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o;
        end else begin
            l_TColl_0_0_1_constprop_o = l_TColl_0_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_0_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o;
        end else begin
            l_TColl_0_0_2_constprop_o = l_TColl_0_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_0_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o;
        end else begin
            l_TColl_0_0_3_constprop_o = l_TColl_0_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_1_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o;
        end else begin
            l_TColl_0_1_0_constprop_o = l_TColl_0_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_1_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o;
        end else begin
            l_TColl_0_1_1_constprop_o = l_TColl_0_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_1_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o;
        end else begin
            l_TColl_0_1_2_constprop_o = l_TColl_0_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_1_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o;
        end else begin
            l_TColl_0_1_3_constprop_o = l_TColl_0_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_2_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o;
        end else begin
            l_TColl_0_2_0_constprop_o = l_TColl_0_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_2_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o;
        end else begin
            l_TColl_0_2_1_constprop_o = l_TColl_0_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_2_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o;
        end else begin
            l_TColl_0_2_2_constprop_o = l_TColl_0_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_2_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o;
        end else begin
            l_TColl_0_2_3_constprop_o = l_TColl_0_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_3_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o;
        end else begin
            l_TColl_0_3_0_constprop_o = l_TColl_0_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_3_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o;
        end else begin
            l_TColl_0_3_1_constprop_o = l_TColl_0_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_3_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o;
        end else begin
            l_TColl_0_3_2_constprop_o = l_TColl_0_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_0_3_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o;
        end else begin
            l_TColl_0_3_3_constprop_o = l_TColl_0_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_0_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o;
        end else begin
            l_TColl_1_0_0_constprop_o = l_TColl_1_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_0_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o;
        end else begin
            l_TColl_1_0_1_constprop_o = l_TColl_1_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_0_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o;
        end else begin
            l_TColl_1_0_2_constprop_o = l_TColl_1_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_0_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o;
        end else begin
            l_TColl_1_0_3_constprop_o = l_TColl_1_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_1_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o;
        end else begin
            l_TColl_1_1_0_constprop_o = l_TColl_1_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_1_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o;
        end else begin
            l_TColl_1_1_1_constprop_o = l_TColl_1_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_1_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o;
        end else begin
            l_TColl_1_1_2_constprop_o = l_TColl_1_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_1_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o;
        end else begin
            l_TColl_1_1_3_constprop_o = l_TColl_1_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_2_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o;
        end else begin
            l_TColl_1_2_0_constprop_o = l_TColl_1_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_2_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o;
        end else begin
            l_TColl_1_2_1_constprop_o = l_TColl_1_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_2_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o;
        end else begin
            l_TColl_1_2_2_constprop_o = l_TColl_1_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_2_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o;
        end else begin
            l_TColl_1_2_3_constprop_o = l_TColl_1_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_3_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o;
        end else begin
            l_TColl_1_3_0_constprop_o = l_TColl_1_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_3_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o;
        end else begin
            l_TColl_1_3_1_constprop_o = l_TColl_1_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_3_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o;
        end else begin
            l_TColl_1_3_2_constprop_o = l_TColl_1_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_1_3_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o;
        end else begin
            l_TColl_1_3_3_constprop_o = l_TColl_1_3_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_0_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o;
        end else begin
            l_TColl_2_0_0_constprop_o = l_TColl_2_0_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_0_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o;
        end else begin
            l_TColl_2_0_1_constprop_o = l_TColl_2_0_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_0_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o;
        end else begin
            l_TColl_2_0_2_constprop_o = l_TColl_2_0_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_0_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o;
        end else begin
            l_TColl_2_0_3_constprop_o = l_TColl_2_0_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_1_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o;
        end else begin
            l_TColl_2_1_0_constprop_o = l_TColl_2_1_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_1_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o;
        end else begin
            l_TColl_2_1_1_constprop_o = l_TColl_2_1_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_1_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o;
        end else begin
            l_TColl_2_1_2_constprop_o = l_TColl_2_1_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_1_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o;
        end else begin
            l_TColl_2_1_3_constprop_o = l_TColl_2_1_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_2_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o;
        end else begin
            l_TColl_2_2_0_constprop_o = l_TColl_2_2_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_2_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o;
        end else begin
            l_TColl_2_2_1_constprop_o = l_TColl_2_2_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_2_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o;
        end else begin
            l_TColl_2_2_2_constprop_o = l_TColl_2_2_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_2_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o;
        end else begin
            l_TColl_2_2_3_constprop_o = l_TColl_2_2_3_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_3_0_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o;
        end else begin
            l_TColl_2_3_0_constprop_o = l_TColl_2_3_0_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_3_1_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o;
        end else begin
            l_TColl_2_3_1_constprop_o = l_TColl_2_3_1_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_3_2_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o;
        end else begin
            l_TColl_2_3_2_constprop_o = l_TColl_2_3_2_constprop_i;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state209))) begin
            l_TColl_2_3_3_constprop_o = grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o;
        end else begin
            l_TColl_2_3_3_constprop_o = l_TColl_2_3_3_constprop_i;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state216)) begin
            qConnect_address0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_address0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            qConnect_address0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_address0;
        end else if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qConnect_address0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_address0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qConnect_address0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_address0;
        end else begin
            qConnect_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state216)) begin
            qConnect_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_qConnect_ce0;
        end else if ((1'b1 == ap_CS_fsm_state207)) begin
            qConnect_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qConnect_ce0;
        end else if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qConnect_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_ce0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qConnect_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_ce0;
        end else begin
            qConnect_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qConnect_d0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_d0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qConnect_d0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_d0;
        end else begin
            qConnect_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qConnect_we0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qConnect_we0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qConnect_we0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qConnect_we0;
        end else begin
            qConnect_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state207)) begin
            qNear_address0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_address0;
        end else if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qNear_address0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_address0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            qNear_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_address0;
        end else if ((1'b1 == ap_CS_fsm_state83)) begin
            qNear_address0 = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_address0;
        end else begin
            qNear_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state207)) begin
            qNear_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_qNear_ce0;
        end else if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qNear_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qNear_ce0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            qNear_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qNear_ce0;
        end else if ((1'b1 == ap_CS_fsm_state83)) begin
            qNear_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_ce0;
        end else begin
            qNear_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state83)) begin
            qNear_we0 = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_qNear_we0;
        end else begin
            qNear_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_address0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_address0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_address0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_address0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_address0;
        end else if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_address0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            qRand_address0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_address0;
        end else begin
            qRand_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln119_reg_2458) & (1'b1 == ap_CS_fsm_state204))) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_qRand_ce0;
        end else if ((1'b1 == ap_CS_fsm_state145)) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_qRand_ce0;
        end else if ((1'b1 == ap_CS_fsm_state85)) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_qRand_ce0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_qRand_ce0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_qRand_ce0;
        end else if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_ce0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            qRand_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_ce0;
        end else begin
            qRand_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            qRand_d0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_d0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            qRand_d0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_d0;
        end else begin
            qRand_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'd1 == and_ln110_reg_2427) & (1'b1 == ap_CS_fsm_state20))) begin
            qRand_we0 = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_qRand_we0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            qRand_we0 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_qRand_we0;
        end else begin
            qRand_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state278)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state216)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state83)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            rrtVertices_address0 = grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_address0;
        end else begin
            rrtVertices_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state278)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state276)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state217)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state216)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state83)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state81)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state22)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_rrtVertices_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            rrtVertices_ce0 = grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_ce0;
        end else begin
            rrtVertices_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            rrtVertices_d0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_d0;
        end else if ((1'b1 == ap_CS_fsm_state216)) begin
            rrtVertices_d0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_d0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            rrtVertices_d0 = grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_d0;
        end else begin
            rrtVertices_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state338) & (icmp_ln107_reg_2379 == 1'd1))) begin
            rrtVertices_we0 = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_rrtVertices_we0;
        end else if ((1'b1 == ap_CS_fsm_state216)) begin
            rrtVertices_we0 = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_rrtVertices_we0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            rrtVertices_we0 = grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_rrtVertices_we0;
        end else begin
            rrtVertices_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                if (((1'b1 == ap_CS_fsm_state2) & (grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end
            end
            ap_ST_fsm_state3: begin
                if (((1'b1 == ap_CS_fsm_state3) & (icmp_ln107_fu_1491_p2 == 1'd0))) begin
                    ap_NS_fsm = ap_ST_fsm_state338;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            ap_ST_fsm_state4: begin
                if (((1'b1 == ap_CS_fsm_state4) & (grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                if (((1'b0 == ap_block_state20_on_subcall_done) & (1'b1 == ap_CS_fsm_state20))) begin
                    ap_NS_fsm = ap_ST_fsm_state21;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state20;
                end
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                if (((1'b1 == ap_CS_fsm_state22) & (grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state23;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state22;
                end
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end
            ap_ST_fsm_state78: begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
            ap_ST_fsm_state79: begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end
            ap_ST_fsm_state80: begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
            ap_ST_fsm_state81: begin
                if (((1'b1 == ap_CS_fsm_state81) & (grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state82;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state81;
                end
            end
            ap_ST_fsm_state82: begin
                ap_NS_fsm = ap_ST_fsm_state83;
            end
            ap_ST_fsm_state83: begin
                if (((1'b1 == ap_CS_fsm_state83) & (grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state84;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state83;
                end
            end
            ap_ST_fsm_state84: begin
                ap_NS_fsm = ap_ST_fsm_state85;
            end
            ap_ST_fsm_state85: begin
                if (((1'b1 == ap_CS_fsm_state85) & (grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state86;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state85;
                end
            end
            ap_ST_fsm_state86: begin
                ap_NS_fsm = ap_ST_fsm_state87;
            end
            ap_ST_fsm_state87: begin
                ap_NS_fsm = ap_ST_fsm_state88;
            end
            ap_ST_fsm_state88: begin
                ap_NS_fsm = ap_ST_fsm_state89;
            end
            ap_ST_fsm_state89: begin
                ap_NS_fsm = ap_ST_fsm_state90;
            end
            ap_ST_fsm_state90: begin
                ap_NS_fsm = ap_ST_fsm_state91;
            end
            ap_ST_fsm_state91: begin
                ap_NS_fsm = ap_ST_fsm_state92;
            end
            ap_ST_fsm_state92: begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end
            ap_ST_fsm_state93: begin
                ap_NS_fsm = ap_ST_fsm_state94;
            end
            ap_ST_fsm_state94: begin
                ap_NS_fsm = ap_ST_fsm_state95;
            end
            ap_ST_fsm_state95: begin
                ap_NS_fsm = ap_ST_fsm_state96;
            end
            ap_ST_fsm_state96: begin
                ap_NS_fsm = ap_ST_fsm_state97;
            end
            ap_ST_fsm_state97: begin
                ap_NS_fsm = ap_ST_fsm_state98;
            end
            ap_ST_fsm_state98: begin
                ap_NS_fsm = ap_ST_fsm_state99;
            end
            ap_ST_fsm_state99: begin
                ap_NS_fsm = ap_ST_fsm_state100;
            end
            ap_ST_fsm_state100: begin
                ap_NS_fsm = ap_ST_fsm_state101;
            end
            ap_ST_fsm_state101: begin
                ap_NS_fsm = ap_ST_fsm_state102;
            end
            ap_ST_fsm_state102: begin
                ap_NS_fsm = ap_ST_fsm_state103;
            end
            ap_ST_fsm_state103: begin
                ap_NS_fsm = ap_ST_fsm_state104;
            end
            ap_ST_fsm_state104: begin
                ap_NS_fsm = ap_ST_fsm_state105;
            end
            ap_ST_fsm_state105: begin
                ap_NS_fsm = ap_ST_fsm_state106;
            end
            ap_ST_fsm_state106: begin
                ap_NS_fsm = ap_ST_fsm_state107;
            end
            ap_ST_fsm_state107: begin
                ap_NS_fsm = ap_ST_fsm_state108;
            end
            ap_ST_fsm_state108: begin
                ap_NS_fsm = ap_ST_fsm_state109;
            end
            ap_ST_fsm_state109: begin
                ap_NS_fsm = ap_ST_fsm_state110;
            end
            ap_ST_fsm_state110: begin
                ap_NS_fsm = ap_ST_fsm_state111;
            end
            ap_ST_fsm_state111: begin
                ap_NS_fsm = ap_ST_fsm_state112;
            end
            ap_ST_fsm_state112: begin
                ap_NS_fsm = ap_ST_fsm_state113;
            end
            ap_ST_fsm_state113: begin
                ap_NS_fsm = ap_ST_fsm_state114;
            end
            ap_ST_fsm_state114: begin
                ap_NS_fsm = ap_ST_fsm_state115;
            end
            ap_ST_fsm_state115: begin
                ap_NS_fsm = ap_ST_fsm_state116;
            end
            ap_ST_fsm_state116: begin
                ap_NS_fsm = ap_ST_fsm_state117;
            end
            ap_ST_fsm_state117: begin
                ap_NS_fsm = ap_ST_fsm_state118;
            end
            ap_ST_fsm_state118: begin
                ap_NS_fsm = ap_ST_fsm_state119;
            end
            ap_ST_fsm_state119: begin
                ap_NS_fsm = ap_ST_fsm_state120;
            end
            ap_ST_fsm_state120: begin
                ap_NS_fsm = ap_ST_fsm_state121;
            end
            ap_ST_fsm_state121: begin
                ap_NS_fsm = ap_ST_fsm_state122;
            end
            ap_ST_fsm_state122: begin
                ap_NS_fsm = ap_ST_fsm_state123;
            end
            ap_ST_fsm_state123: begin
                ap_NS_fsm = ap_ST_fsm_state124;
            end
            ap_ST_fsm_state124: begin
                ap_NS_fsm = ap_ST_fsm_state125;
            end
            ap_ST_fsm_state125: begin
                ap_NS_fsm = ap_ST_fsm_state126;
            end
            ap_ST_fsm_state126: begin
                ap_NS_fsm = ap_ST_fsm_state127;
            end
            ap_ST_fsm_state127: begin
                ap_NS_fsm = ap_ST_fsm_state128;
            end
            ap_ST_fsm_state128: begin
                ap_NS_fsm = ap_ST_fsm_state129;
            end
            ap_ST_fsm_state129: begin
                ap_NS_fsm = ap_ST_fsm_state130;
            end
            ap_ST_fsm_state130: begin
                ap_NS_fsm = ap_ST_fsm_state131;
            end
            ap_ST_fsm_state131: begin
                ap_NS_fsm = ap_ST_fsm_state132;
            end
            ap_ST_fsm_state132: begin
                ap_NS_fsm = ap_ST_fsm_state133;
            end
            ap_ST_fsm_state133: begin
                ap_NS_fsm = ap_ST_fsm_state134;
            end
            ap_ST_fsm_state134: begin
                ap_NS_fsm = ap_ST_fsm_state135;
            end
            ap_ST_fsm_state135: begin
                ap_NS_fsm = ap_ST_fsm_state136;
            end
            ap_ST_fsm_state136: begin
                ap_NS_fsm = ap_ST_fsm_state137;
            end
            ap_ST_fsm_state137: begin
                ap_NS_fsm = ap_ST_fsm_state138;
            end
            ap_ST_fsm_state138: begin
                ap_NS_fsm = ap_ST_fsm_state139;
            end
            ap_ST_fsm_state139: begin
                ap_NS_fsm = ap_ST_fsm_state140;
            end
            ap_ST_fsm_state140: begin
                ap_NS_fsm = ap_ST_fsm_state141;
            end
            ap_ST_fsm_state141: begin
                ap_NS_fsm = ap_ST_fsm_state142;
            end
            ap_ST_fsm_state142: begin
                ap_NS_fsm = ap_ST_fsm_state143;
            end
            ap_ST_fsm_state143: begin
                ap_NS_fsm = ap_ST_fsm_state144;
            end
            ap_ST_fsm_state144: begin
                if (((1'd1 == and_ln119_fu_1767_p2) & (1'b1 == ap_CS_fsm_state144))) begin
                    ap_NS_fsm = ap_ST_fsm_state146;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state145;
                end
            end
            ap_ST_fsm_state145: begin
                if (((1'b1 == ap_CS_fsm_state145) & (grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state204;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state145;
                end
            end
            ap_ST_fsm_state146: begin
                ap_NS_fsm = ap_ST_fsm_state147;
            end
            ap_ST_fsm_state147: begin
                ap_NS_fsm = ap_ST_fsm_state148;
            end
            ap_ST_fsm_state148: begin
                ap_NS_fsm = ap_ST_fsm_state149;
            end
            ap_ST_fsm_state149: begin
                ap_NS_fsm = ap_ST_fsm_state150;
            end
            ap_ST_fsm_state150: begin
                ap_NS_fsm = ap_ST_fsm_state151;
            end
            ap_ST_fsm_state151: begin
                ap_NS_fsm = ap_ST_fsm_state152;
            end
            ap_ST_fsm_state152: begin
                ap_NS_fsm = ap_ST_fsm_state153;
            end
            ap_ST_fsm_state153: begin
                ap_NS_fsm = ap_ST_fsm_state154;
            end
            ap_ST_fsm_state154: begin
                ap_NS_fsm = ap_ST_fsm_state155;
            end
            ap_ST_fsm_state155: begin
                ap_NS_fsm = ap_ST_fsm_state156;
            end
            ap_ST_fsm_state156: begin
                ap_NS_fsm = ap_ST_fsm_state157;
            end
            ap_ST_fsm_state157: begin
                ap_NS_fsm = ap_ST_fsm_state158;
            end
            ap_ST_fsm_state158: begin
                ap_NS_fsm = ap_ST_fsm_state159;
            end
            ap_ST_fsm_state159: begin
                ap_NS_fsm = ap_ST_fsm_state160;
            end
            ap_ST_fsm_state160: begin
                ap_NS_fsm = ap_ST_fsm_state161;
            end
            ap_ST_fsm_state161: begin
                ap_NS_fsm = ap_ST_fsm_state162;
            end
            ap_ST_fsm_state162: begin
                ap_NS_fsm = ap_ST_fsm_state163;
            end
            ap_ST_fsm_state163: begin
                ap_NS_fsm = ap_ST_fsm_state164;
            end
            ap_ST_fsm_state164: begin
                ap_NS_fsm = ap_ST_fsm_state165;
            end
            ap_ST_fsm_state165: begin
                ap_NS_fsm = ap_ST_fsm_state166;
            end
            ap_ST_fsm_state166: begin
                ap_NS_fsm = ap_ST_fsm_state167;
            end
            ap_ST_fsm_state167: begin
                ap_NS_fsm = ap_ST_fsm_state168;
            end
            ap_ST_fsm_state168: begin
                ap_NS_fsm = ap_ST_fsm_state169;
            end
            ap_ST_fsm_state169: begin
                ap_NS_fsm = ap_ST_fsm_state170;
            end
            ap_ST_fsm_state170: begin
                ap_NS_fsm = ap_ST_fsm_state171;
            end
            ap_ST_fsm_state171: begin
                ap_NS_fsm = ap_ST_fsm_state172;
            end
            ap_ST_fsm_state172: begin
                ap_NS_fsm = ap_ST_fsm_state173;
            end
            ap_ST_fsm_state173: begin
                ap_NS_fsm = ap_ST_fsm_state174;
            end
            ap_ST_fsm_state174: begin
                ap_NS_fsm = ap_ST_fsm_state175;
            end
            ap_ST_fsm_state175: begin
                ap_NS_fsm = ap_ST_fsm_state176;
            end
            ap_ST_fsm_state176: begin
                ap_NS_fsm = ap_ST_fsm_state177;
            end
            ap_ST_fsm_state177: begin
                ap_NS_fsm = ap_ST_fsm_state178;
            end
            ap_ST_fsm_state178: begin
                ap_NS_fsm = ap_ST_fsm_state179;
            end
            ap_ST_fsm_state179: begin
                ap_NS_fsm = ap_ST_fsm_state180;
            end
            ap_ST_fsm_state180: begin
                ap_NS_fsm = ap_ST_fsm_state181;
            end
            ap_ST_fsm_state181: begin
                ap_NS_fsm = ap_ST_fsm_state182;
            end
            ap_ST_fsm_state182: begin
                ap_NS_fsm = ap_ST_fsm_state183;
            end
            ap_ST_fsm_state183: begin
                ap_NS_fsm = ap_ST_fsm_state184;
            end
            ap_ST_fsm_state184: begin
                ap_NS_fsm = ap_ST_fsm_state185;
            end
            ap_ST_fsm_state185: begin
                ap_NS_fsm = ap_ST_fsm_state186;
            end
            ap_ST_fsm_state186: begin
                ap_NS_fsm = ap_ST_fsm_state187;
            end
            ap_ST_fsm_state187: begin
                ap_NS_fsm = ap_ST_fsm_state188;
            end
            ap_ST_fsm_state188: begin
                ap_NS_fsm = ap_ST_fsm_state189;
            end
            ap_ST_fsm_state189: begin
                ap_NS_fsm = ap_ST_fsm_state190;
            end
            ap_ST_fsm_state190: begin
                ap_NS_fsm = ap_ST_fsm_state191;
            end
            ap_ST_fsm_state191: begin
                ap_NS_fsm = ap_ST_fsm_state192;
            end
            ap_ST_fsm_state192: begin
                ap_NS_fsm = ap_ST_fsm_state193;
            end
            ap_ST_fsm_state193: begin
                ap_NS_fsm = ap_ST_fsm_state194;
            end
            ap_ST_fsm_state194: begin
                ap_NS_fsm = ap_ST_fsm_state195;
            end
            ap_ST_fsm_state195: begin
                ap_NS_fsm = ap_ST_fsm_state196;
            end
            ap_ST_fsm_state196: begin
                ap_NS_fsm = ap_ST_fsm_state197;
            end
            ap_ST_fsm_state197: begin
                ap_NS_fsm = ap_ST_fsm_state198;
            end
            ap_ST_fsm_state198: begin
                ap_NS_fsm = ap_ST_fsm_state199;
            end
            ap_ST_fsm_state199: begin
                ap_NS_fsm = ap_ST_fsm_state200;
            end
            ap_ST_fsm_state200: begin
                ap_NS_fsm = ap_ST_fsm_state201;
            end
            ap_ST_fsm_state201: begin
                ap_NS_fsm = ap_ST_fsm_state202;
            end
            ap_ST_fsm_state202: begin
                ap_NS_fsm = ap_ST_fsm_state203;
            end
            ap_ST_fsm_state203: begin
                ap_NS_fsm = ap_ST_fsm_state204;
            end
            ap_ST_fsm_state204: begin
                if (((1'b0 == ap_block_state204_on_subcall_done) & (1'b1 == ap_CS_fsm_state204))) begin
                    ap_NS_fsm = ap_ST_fsm_state205;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state204;
                end
            end
            ap_ST_fsm_state205: begin
                ap_NS_fsm = ap_ST_fsm_state206;
            end
            ap_ST_fsm_state206: begin
                if (((1'd0 == and_ln188_fu_1809_p2) & (1'b1 == ap_CS_fsm_state206))) begin
                    ap_NS_fsm = ap_ST_fsm_state216;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state207;
                end
            end
            ap_ST_fsm_state207: begin
                if (((1'b1 == ap_CS_fsm_state207) & (grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state208;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state207;
                end
            end
            ap_ST_fsm_state208: begin
                ap_NS_fsm = ap_ST_fsm_state209;
            end
            ap_ST_fsm_state209: begin
                if (((1'b0 == ap_block_state209_on_subcall_done) & (1'b1 == ap_CS_fsm_state209) & ((1'd0 == and_ln188_reg_2467) | (grp_detectCollNode_fu_1055_ap_return == 1'd1)))) begin
                    ap_NS_fsm = ap_ST_fsm_state217;
                end else if (((1'b0 == ap_block_state209_on_subcall_done) & (1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state209))) begin
                    ap_NS_fsm = ap_ST_fsm_state210;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state209;
                end
            end
            ap_ST_fsm_state210: begin
                ap_NS_fsm = ap_ST_fsm_state211;
            end
            ap_ST_fsm_state211: begin
                ap_NS_fsm = ap_ST_fsm_state212;
            end
            ap_ST_fsm_state212: begin
                ap_NS_fsm = ap_ST_fsm_state213;
            end
            ap_ST_fsm_state213: begin
                ap_NS_fsm = ap_ST_fsm_state214;
            end
            ap_ST_fsm_state214: begin
                ap_NS_fsm = ap_ST_fsm_state215;
            end
            ap_ST_fsm_state215: begin
                ap_NS_fsm = ap_ST_fsm_state205;
            end
            ap_ST_fsm_state216: begin
                if (((1'b1 == ap_CS_fsm_state216) & (grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state209;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state216;
                end
            end
            ap_ST_fsm_state217: begin
                if (((grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state217))) begin
                    ap_NS_fsm = ap_ST_fsm_state218;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state217;
                end
            end
            ap_ST_fsm_state218: begin
                ap_NS_fsm = ap_ST_fsm_state219;
            end
            ap_ST_fsm_state219: begin
                ap_NS_fsm = ap_ST_fsm_state220;
            end
            ap_ST_fsm_state220: begin
                ap_NS_fsm = ap_ST_fsm_state221;
            end
            ap_ST_fsm_state221: begin
                ap_NS_fsm = ap_ST_fsm_state222;
            end
            ap_ST_fsm_state222: begin
                ap_NS_fsm = ap_ST_fsm_state223;
            end
            ap_ST_fsm_state223: begin
                ap_NS_fsm = ap_ST_fsm_state224;
            end
            ap_ST_fsm_state224: begin
                ap_NS_fsm = ap_ST_fsm_state225;
            end
            ap_ST_fsm_state225: begin
                ap_NS_fsm = ap_ST_fsm_state226;
            end
            ap_ST_fsm_state226: begin
                ap_NS_fsm = ap_ST_fsm_state227;
            end
            ap_ST_fsm_state227: begin
                ap_NS_fsm = ap_ST_fsm_state228;
            end
            ap_ST_fsm_state228: begin
                ap_NS_fsm = ap_ST_fsm_state229;
            end
            ap_ST_fsm_state229: begin
                ap_NS_fsm = ap_ST_fsm_state230;
            end
            ap_ST_fsm_state230: begin
                ap_NS_fsm = ap_ST_fsm_state231;
            end
            ap_ST_fsm_state231: begin
                ap_NS_fsm = ap_ST_fsm_state232;
            end
            ap_ST_fsm_state232: begin
                ap_NS_fsm = ap_ST_fsm_state233;
            end
            ap_ST_fsm_state233: begin
                ap_NS_fsm = ap_ST_fsm_state234;
            end
            ap_ST_fsm_state234: begin
                ap_NS_fsm = ap_ST_fsm_state235;
            end
            ap_ST_fsm_state235: begin
                ap_NS_fsm = ap_ST_fsm_state236;
            end
            ap_ST_fsm_state236: begin
                ap_NS_fsm = ap_ST_fsm_state237;
            end
            ap_ST_fsm_state237: begin
                ap_NS_fsm = ap_ST_fsm_state238;
            end
            ap_ST_fsm_state238: begin
                ap_NS_fsm = ap_ST_fsm_state239;
            end
            ap_ST_fsm_state239: begin
                ap_NS_fsm = ap_ST_fsm_state240;
            end
            ap_ST_fsm_state240: begin
                ap_NS_fsm = ap_ST_fsm_state241;
            end
            ap_ST_fsm_state241: begin
                ap_NS_fsm = ap_ST_fsm_state242;
            end
            ap_ST_fsm_state242: begin
                ap_NS_fsm = ap_ST_fsm_state243;
            end
            ap_ST_fsm_state243: begin
                ap_NS_fsm = ap_ST_fsm_state244;
            end
            ap_ST_fsm_state244: begin
                ap_NS_fsm = ap_ST_fsm_state245;
            end
            ap_ST_fsm_state245: begin
                ap_NS_fsm = ap_ST_fsm_state246;
            end
            ap_ST_fsm_state246: begin
                ap_NS_fsm = ap_ST_fsm_state247;
            end
            ap_ST_fsm_state247: begin
                ap_NS_fsm = ap_ST_fsm_state248;
            end
            ap_ST_fsm_state248: begin
                ap_NS_fsm = ap_ST_fsm_state249;
            end
            ap_ST_fsm_state249: begin
                ap_NS_fsm = ap_ST_fsm_state250;
            end
            ap_ST_fsm_state250: begin
                ap_NS_fsm = ap_ST_fsm_state251;
            end
            ap_ST_fsm_state251: begin
                ap_NS_fsm = ap_ST_fsm_state252;
            end
            ap_ST_fsm_state252: begin
                ap_NS_fsm = ap_ST_fsm_state253;
            end
            ap_ST_fsm_state253: begin
                ap_NS_fsm = ap_ST_fsm_state254;
            end
            ap_ST_fsm_state254: begin
                ap_NS_fsm = ap_ST_fsm_state255;
            end
            ap_ST_fsm_state255: begin
                ap_NS_fsm = ap_ST_fsm_state256;
            end
            ap_ST_fsm_state256: begin
                ap_NS_fsm = ap_ST_fsm_state257;
            end
            ap_ST_fsm_state257: begin
                ap_NS_fsm = ap_ST_fsm_state258;
            end
            ap_ST_fsm_state258: begin
                ap_NS_fsm = ap_ST_fsm_state259;
            end
            ap_ST_fsm_state259: begin
                ap_NS_fsm = ap_ST_fsm_state260;
            end
            ap_ST_fsm_state260: begin
                ap_NS_fsm = ap_ST_fsm_state261;
            end
            ap_ST_fsm_state261: begin
                ap_NS_fsm = ap_ST_fsm_state262;
            end
            ap_ST_fsm_state262: begin
                ap_NS_fsm = ap_ST_fsm_state263;
            end
            ap_ST_fsm_state263: begin
                ap_NS_fsm = ap_ST_fsm_state264;
            end
            ap_ST_fsm_state264: begin
                ap_NS_fsm = ap_ST_fsm_state265;
            end
            ap_ST_fsm_state265: begin
                ap_NS_fsm = ap_ST_fsm_state266;
            end
            ap_ST_fsm_state266: begin
                ap_NS_fsm = ap_ST_fsm_state267;
            end
            ap_ST_fsm_state267: begin
                ap_NS_fsm = ap_ST_fsm_state268;
            end
            ap_ST_fsm_state268: begin
                ap_NS_fsm = ap_ST_fsm_state269;
            end
            ap_ST_fsm_state269: begin
                ap_NS_fsm = ap_ST_fsm_state270;
            end
            ap_ST_fsm_state270: begin
                ap_NS_fsm = ap_ST_fsm_state271;
            end
            ap_ST_fsm_state271: begin
                ap_NS_fsm = ap_ST_fsm_state272;
            end
            ap_ST_fsm_state272: begin
                ap_NS_fsm = ap_ST_fsm_state273;
            end
            ap_ST_fsm_state273: begin
                ap_NS_fsm = ap_ST_fsm_state274;
            end
            ap_ST_fsm_state274: begin
                ap_NS_fsm = ap_ST_fsm_state275;
            end
            ap_ST_fsm_state275: begin
                ap_NS_fsm = ap_ST_fsm_state276;
            end
            ap_ST_fsm_state276: begin
                if (((grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state276))) begin
                    ap_NS_fsm = ap_ST_fsm_state277;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state276;
                end
            end
            ap_ST_fsm_state277: begin
                ap_NS_fsm = ap_ST_fsm_state278;
            end
            ap_ST_fsm_state278: begin
                if (((grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state278))) begin
                    ap_NS_fsm = ap_ST_fsm_state279;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state278;
                end
            end
            ap_ST_fsm_state279: begin
                ap_NS_fsm = ap_ST_fsm_state280;
            end
            ap_ST_fsm_state280: begin
                ap_NS_fsm = ap_ST_fsm_state281;
            end
            ap_ST_fsm_state281: begin
                ap_NS_fsm = ap_ST_fsm_state282;
            end
            ap_ST_fsm_state282: begin
                ap_NS_fsm = ap_ST_fsm_state283;
            end
            ap_ST_fsm_state283: begin
                ap_NS_fsm = ap_ST_fsm_state284;
            end
            ap_ST_fsm_state284: begin
                ap_NS_fsm = ap_ST_fsm_state285;
            end
            ap_ST_fsm_state285: begin
                ap_NS_fsm = ap_ST_fsm_state286;
            end
            ap_ST_fsm_state286: begin
                ap_NS_fsm = ap_ST_fsm_state287;
            end
            ap_ST_fsm_state287: begin
                ap_NS_fsm = ap_ST_fsm_state288;
            end
            ap_ST_fsm_state288: begin
                ap_NS_fsm = ap_ST_fsm_state289;
            end
            ap_ST_fsm_state289: begin
                ap_NS_fsm = ap_ST_fsm_state290;
            end
            ap_ST_fsm_state290: begin
                ap_NS_fsm = ap_ST_fsm_state291;
            end
            ap_ST_fsm_state291: begin
                ap_NS_fsm = ap_ST_fsm_state292;
            end
            ap_ST_fsm_state292: begin
                ap_NS_fsm = ap_ST_fsm_state293;
            end
            ap_ST_fsm_state293: begin
                ap_NS_fsm = ap_ST_fsm_state294;
            end
            ap_ST_fsm_state294: begin
                ap_NS_fsm = ap_ST_fsm_state295;
            end
            ap_ST_fsm_state295: begin
                ap_NS_fsm = ap_ST_fsm_state296;
            end
            ap_ST_fsm_state296: begin
                ap_NS_fsm = ap_ST_fsm_state297;
            end
            ap_ST_fsm_state297: begin
                ap_NS_fsm = ap_ST_fsm_state298;
            end
            ap_ST_fsm_state298: begin
                ap_NS_fsm = ap_ST_fsm_state299;
            end
            ap_ST_fsm_state299: begin
                ap_NS_fsm = ap_ST_fsm_state300;
            end
            ap_ST_fsm_state300: begin
                ap_NS_fsm = ap_ST_fsm_state301;
            end
            ap_ST_fsm_state301: begin
                ap_NS_fsm = ap_ST_fsm_state302;
            end
            ap_ST_fsm_state302: begin
                ap_NS_fsm = ap_ST_fsm_state303;
            end
            ap_ST_fsm_state303: begin
                ap_NS_fsm = ap_ST_fsm_state304;
            end
            ap_ST_fsm_state304: begin
                ap_NS_fsm = ap_ST_fsm_state305;
            end
            ap_ST_fsm_state305: begin
                ap_NS_fsm = ap_ST_fsm_state306;
            end
            ap_ST_fsm_state306: begin
                ap_NS_fsm = ap_ST_fsm_state307;
            end
            ap_ST_fsm_state307: begin
                ap_NS_fsm = ap_ST_fsm_state308;
            end
            ap_ST_fsm_state308: begin
                ap_NS_fsm = ap_ST_fsm_state309;
            end
            ap_ST_fsm_state309: begin
                ap_NS_fsm = ap_ST_fsm_state310;
            end
            ap_ST_fsm_state310: begin
                ap_NS_fsm = ap_ST_fsm_state311;
            end
            ap_ST_fsm_state311: begin
                ap_NS_fsm = ap_ST_fsm_state312;
            end
            ap_ST_fsm_state312: begin
                ap_NS_fsm = ap_ST_fsm_state313;
            end
            ap_ST_fsm_state313: begin
                ap_NS_fsm = ap_ST_fsm_state314;
            end
            ap_ST_fsm_state314: begin
                ap_NS_fsm = ap_ST_fsm_state315;
            end
            ap_ST_fsm_state315: begin
                ap_NS_fsm = ap_ST_fsm_state316;
            end
            ap_ST_fsm_state316: begin
                ap_NS_fsm = ap_ST_fsm_state317;
            end
            ap_ST_fsm_state317: begin
                ap_NS_fsm = ap_ST_fsm_state318;
            end
            ap_ST_fsm_state318: begin
                ap_NS_fsm = ap_ST_fsm_state319;
            end
            ap_ST_fsm_state319: begin
                ap_NS_fsm = ap_ST_fsm_state320;
            end
            ap_ST_fsm_state320: begin
                ap_NS_fsm = ap_ST_fsm_state321;
            end
            ap_ST_fsm_state321: begin
                ap_NS_fsm = ap_ST_fsm_state322;
            end
            ap_ST_fsm_state322: begin
                ap_NS_fsm = ap_ST_fsm_state323;
            end
            ap_ST_fsm_state323: begin
                ap_NS_fsm = ap_ST_fsm_state324;
            end
            ap_ST_fsm_state324: begin
                ap_NS_fsm = ap_ST_fsm_state325;
            end
            ap_ST_fsm_state325: begin
                ap_NS_fsm = ap_ST_fsm_state326;
            end
            ap_ST_fsm_state326: begin
                ap_NS_fsm = ap_ST_fsm_state327;
            end
            ap_ST_fsm_state327: begin
                ap_NS_fsm = ap_ST_fsm_state328;
            end
            ap_ST_fsm_state328: begin
                ap_NS_fsm = ap_ST_fsm_state329;
            end
            ap_ST_fsm_state329: begin
                ap_NS_fsm = ap_ST_fsm_state330;
            end
            ap_ST_fsm_state330: begin
                ap_NS_fsm = ap_ST_fsm_state331;
            end
            ap_ST_fsm_state331: begin
                ap_NS_fsm = ap_ST_fsm_state332;
            end
            ap_ST_fsm_state332: begin
                ap_NS_fsm = ap_ST_fsm_state333;
            end
            ap_ST_fsm_state333: begin
                ap_NS_fsm = ap_ST_fsm_state334;
            end
            ap_ST_fsm_state334: begin
                ap_NS_fsm = ap_ST_fsm_state335;
            end
            ap_ST_fsm_state335: begin
                ap_NS_fsm = ap_ST_fsm_state336;
            end
            ap_ST_fsm_state336: begin
                ap_NS_fsm = ap_ST_fsm_state337;
            end
            ap_ST_fsm_state337: begin
                if (((1'd0 == and_ln138_fu_1960_p2) & (1'b1 == ap_CS_fsm_state337))) begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state338;
                end
            end
            ap_ST_fsm_state338: begin
                if (((1'b0 == ap_block_state338_on_subcall_done) & (1'b1 == ap_CS_fsm_state338))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state338;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln96_2_fu_1659_p2 = ($signed(numVertices_1_reg_2362) + $signed(32'd4294967295));

    assign add_ln96_fu_1853_p2 = ($signed(numVertices_fu_520) + $signed(32'd4294967295));

    assign and_ln110_fu_1614_p2 = (or_ln110_fu_1610_p2 & grp_fu_1454_p2);

    assign and_ln119_fu_1767_p2 = (or_ln119_fu_1761_p2 & grp_fu_1454_p2);

    assign and_ln138_fu_1960_p2 = (or_ln138_fu_1956_p2 & grp_fu_1454_p2);

    assign and_ln188_fu_1809_p2 = (or_ln188_fu_1803_p2 & grp_fu_1454_p2);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state142 = ap_CS_fsm[32'd141];

    assign ap_CS_fsm_state143 = ap_CS_fsm[32'd142];

    assign ap_CS_fsm_state144 = ap_CS_fsm[32'd143];

    assign ap_CS_fsm_state145 = ap_CS_fsm[32'd144];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

    assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

    assign ap_CS_fsm_state203 = ap_CS_fsm[32'd202];

    assign ap_CS_fsm_state204 = ap_CS_fsm[32'd203];

    assign ap_CS_fsm_state205 = ap_CS_fsm[32'd204];

    assign ap_CS_fsm_state206 = ap_CS_fsm[32'd205];

    assign ap_CS_fsm_state207 = ap_CS_fsm[32'd206];

    assign ap_CS_fsm_state208 = ap_CS_fsm[32'd207];

    assign ap_CS_fsm_state209 = ap_CS_fsm[32'd208];

    assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];

    assign ap_CS_fsm_state210 = ap_CS_fsm[32'd209];

    assign ap_CS_fsm_state211 = ap_CS_fsm[32'd210];

    assign ap_CS_fsm_state212 = ap_CS_fsm[32'd211];

    assign ap_CS_fsm_state213 = ap_CS_fsm[32'd212];

    assign ap_CS_fsm_state214 = ap_CS_fsm[32'd213];

    assign ap_CS_fsm_state215 = ap_CS_fsm[32'd214];

    assign ap_CS_fsm_state216 = ap_CS_fsm[32'd215];

    assign ap_CS_fsm_state217 = ap_CS_fsm[32'd216];

    assign ap_CS_fsm_state218 = ap_CS_fsm[32'd217];

    assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];

    assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];

    assign ap_CS_fsm_state274 = ap_CS_fsm[32'd273];

    assign ap_CS_fsm_state275 = ap_CS_fsm[32'd274];

    assign ap_CS_fsm_state276 = ap_CS_fsm[32'd275];

    assign ap_CS_fsm_state277 = ap_CS_fsm[32'd276];

    assign ap_CS_fsm_state278 = ap_CS_fsm[32'd277];

    assign ap_CS_fsm_state279 = ap_CS_fsm[32'd278];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state335 = ap_CS_fsm[32'd334];

    assign ap_CS_fsm_state336 = ap_CS_fsm[32'd335];

    assign ap_CS_fsm_state337 = ap_CS_fsm[32'd336];

    assign ap_CS_fsm_state338 = ap_CS_fsm[32'd337];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

    assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

    assign ap_CS_fsm_state81 = ap_CS_fsm[32'd80];

    assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];

    assign ap_CS_fsm_state83 = ap_CS_fsm[32'd82];

    assign ap_CS_fsm_state84 = ap_CS_fsm[32'd83];

    assign ap_CS_fsm_state85 = ap_CS_fsm[32'd84];

    assign ap_CS_fsm_state86 = ap_CS_fsm[32'd85];

    always @(*) begin
        ap_block_state204_on_subcall_done = ((1'd1 == and_ln119_reg_2458) & (grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_done == 1'b0));
    end

    always @(*) begin
        ap_block_state209_on_subcall_done = ((1'd1 == and_ln188_reg_2467) & (grp_detectCollNode_fu_1055_ap_done == 1'b0));
    end

    always @(*) begin
        ap_block_state20_on_subcall_done = ((1'd1 == and_ln110_reg_2427) & (grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_done == 1'b0));
    end

    always @(*) begin
        ap_block_state338_on_subcall_done = ((grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_done == 1'b0) & (icmp_ln107_reg_2379 == 1'd1));
    end

    assign bitcast_ln110_fu_1581_p1 = conv_reg_2411;

    assign bitcast_ln119_fu_1731_p1 = reg_1470;

    assign bitcast_ln138_fu_1926_p1 = reg_1470;

    assign bitcast_ln188_fu_1773_p1 = s_reg_960;

    assign empty_64_fu_1895_p1 = bestIdx_6_loc_fu_528[9:0];

    assign empty_fu_1700_p1 = bestIdx_3_loc_fu_540[9:0];

    assign grp_detectCollNode_fu_1055_ap_start = grp_detectCollNode_fu_1055_ap_start_reg;

    assign grp_fu_2403_p_ce = grp_fu_2529_ce;

    assign grp_fu_2403_p_din0 = grp_fu_2529_p0;

    assign grp_fu_2403_p_din1 = grp_fu_2529_p1;

    assign grp_fu_2403_p_opcode = grp_fu_2529_opcode;

    assign grp_fu_2407_p_ce = grp_fu_2537_ce;

    assign grp_fu_2407_p_din0 = grp_fu_2537_p0;

    assign grp_fu_2407_p_din1 = grp_fu_2537_p1;

    assign grp_fu_2407_p_opcode = grp_fu_2537_opcode;

    assign grp_fu_2411_p_ce = grp_fu_2541_ce;

    assign grp_fu_2411_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2541_p_din0;

    assign grp_fu_2411_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2541_p_din1;

    assign grp_fu_2411_p_opcode = grp_detectCollNode_fu_1055_grp_fu_2541_p_opcode;

    assign grp_fu_2415_p_ce = grp_fu_2545_ce;

    assign grp_fu_2415_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2545_p_din0;

    assign grp_fu_2415_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2545_p_din1;

    assign grp_fu_2415_p_opcode = 2'd0;

    assign grp_fu_2419_p_ce = grp_fu_2549_ce;

    assign grp_fu_2419_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2549_p_din0;

    assign grp_fu_2419_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2549_p_din1;

    assign grp_fu_2419_p_opcode = 2'd0;

    assign grp_fu_2423_p_ce = grp_fu_2553_ce;

    assign grp_fu_2423_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2553_p_din0;

    assign grp_fu_2423_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2553_p_din1;

    assign grp_fu_2423_p_opcode = 2'd0;

    assign grp_fu_2427_p_ce = grp_fu_1442_ce;

    assign grp_fu_2427_p_din0 = s_reg_960;

    assign grp_fu_2427_p_din1 = 64'd4598175219545276416;

    assign grp_fu_2427_p_opcode = 2'd0;

    assign grp_fu_2431_p_ce = grp_fu_2533_ce;

    assign grp_fu_2431_p_din0 = grp_fu_2533_p0;

    assign grp_fu_2431_p_din1 = grp_fu_2533_p1;

    assign grp_fu_2435_p_ce = grp_fu_2557_ce;

    assign grp_fu_2435_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2557_p_din0;

    assign grp_fu_2435_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2557_p_din1;

    assign grp_fu_2439_p_ce = grp_fu_2561_ce;

    assign grp_fu_2439_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2561_p_din0;

    assign grp_fu_2439_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2561_p_din1;

    assign grp_fu_2443_p_ce = grp_fu_2565_ce;

    assign grp_fu_2443_p_din0 = grp_detectCollNode_fu_1055_grp_fu_2565_p_din0;

    assign grp_fu_2443_p_din1 = grp_detectCollNode_fu_1055_grp_fu_2565_p_din1;

    assign grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_110_4_fu_988_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_114_5_fu_1011_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_121_6_fu_1031_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_125_7_fu_1025_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_130_8_fu_1048_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_139_9_fu_1423_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_190_2_fu_1039_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_293_111_fu_1414_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_293_18_fu_1018_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_293_19_fu_1396_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_293_1_fu_995_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_86_1_fu_972_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110_fu_1404_ap_start_reg;

    assign grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start = grp_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1_fu_1002_ap_start_reg;

    assign icmp35_fu_1847_p2 = (($signed(tmp_20_fu_1837_p4) > $signed(31'd0)) ? 1'b1 : 1'b0);

    assign icmp_fu_1653_p2 = (($signed(tmp_19_fu_1644_p4) > $signed(31'd0)) ? 1'b1 : 1'b0);

    assign icmp_ln107_fu_1491_p2 = (($signed(
        numVertices_fu_520
    ) < $signed(
        32'd3000
    )) ? 1'b1 : 1'b0);

    assign icmp_ln110_1_fu_1604_p2 = ((trunc_ln110_fu_1594_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln110_fu_1598_p2 = ((tmp_262_fu_1584_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln119_1_fu_1755_p2 = ((trunc_ln119_fu_1745_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln119_fu_1749_p2 = ((tmp_264_fu_1735_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln138_1_fu_1950_p2 = ((trunc_ln138_fu_1940_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln138_fu_1944_p2 = ((tmp_268_fu_1930_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln188_1_fu_1797_p2 = ((trunc_ln188_fu_1787_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln188_fu_1791_p2 = ((tmp_266_fu_1777_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign l_TColl_0_0_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_0_0_constprop_o_ap_vld;

    assign l_TColl_0_0_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_0_1_constprop_o_ap_vld;

    assign l_TColl_0_0_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_0_2_constprop_o_ap_vld;

    assign l_TColl_0_0_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_0_3_constprop_o_ap_vld;

    assign l_TColl_0_1_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_1_0_constprop_o_ap_vld;

    assign l_TColl_0_1_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_1_1_constprop_o_ap_vld;

    assign l_TColl_0_1_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_1_2_constprop_o_ap_vld;

    assign l_TColl_0_1_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_1_3_constprop_o_ap_vld;

    assign l_TColl_0_2_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_2_0_constprop_o_ap_vld;

    assign l_TColl_0_2_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_2_1_constprop_o_ap_vld;

    assign l_TColl_0_2_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_2_2_constprop_o_ap_vld;

    assign l_TColl_0_2_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_2_3_constprop_o_ap_vld;

    assign l_TColl_0_3_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_3_0_constprop_o_ap_vld;

    assign l_TColl_0_3_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_3_1_constprop_o_ap_vld;

    assign l_TColl_0_3_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_3_2_constprop_o_ap_vld;

    assign l_TColl_0_3_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_0_3_3_constprop_o_ap_vld;

    assign l_TColl_1_0_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_0_0_constprop_o_ap_vld;

    assign l_TColl_1_0_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_0_1_constprop_o_ap_vld;

    assign l_TColl_1_0_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_0_2_constprop_o_ap_vld;

    assign l_TColl_1_0_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_0_3_constprop_o_ap_vld;

    assign l_TColl_1_1_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_1_0_constprop_o_ap_vld;

    assign l_TColl_1_1_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_1_1_constprop_o_ap_vld;

    assign l_TColl_1_1_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_1_2_constprop_o_ap_vld;

    assign l_TColl_1_1_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_1_3_constprop_o_ap_vld;

    assign l_TColl_1_2_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_2_0_constprop_o_ap_vld;

    assign l_TColl_1_2_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_2_1_constprop_o_ap_vld;

    assign l_TColl_1_2_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_2_2_constprop_o_ap_vld;

    assign l_TColl_1_2_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_2_3_constprop_o_ap_vld;

    assign l_TColl_1_3_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_3_0_constprop_o_ap_vld;

    assign l_TColl_1_3_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_3_1_constprop_o_ap_vld;

    assign l_TColl_1_3_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_3_2_constprop_o_ap_vld;

    assign l_TColl_1_3_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_1_3_3_constprop_o_ap_vld;

    assign l_TColl_2_0_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_0_0_constprop_o_ap_vld;

    assign l_TColl_2_0_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_0_1_constprop_o_ap_vld;

    assign l_TColl_2_0_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_0_2_constprop_o_ap_vld;

    assign l_TColl_2_0_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_0_3_constprop_o_ap_vld;

    assign l_TColl_2_1_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_1_0_constprop_o_ap_vld;

    assign l_TColl_2_1_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_1_1_constprop_o_ap_vld;

    assign l_TColl_2_1_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_1_2_constprop_o_ap_vld;

    assign l_TColl_2_1_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_1_3_constprop_o_ap_vld;

    assign l_TColl_2_2_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_2_0_constprop_o_ap_vld;

    assign l_TColl_2_2_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_2_1_constprop_o_ap_vld;

    assign l_TColl_2_2_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_2_2_constprop_o_ap_vld;

    assign l_TColl_2_2_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_2_3_constprop_o_ap_vld;

    assign l_TColl_2_3_0_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_3_0_constprop_o_ap_vld;

    assign l_TColl_2_3_1_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_3_1_constprop_o_ap_vld;

    assign l_TColl_2_3_2_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_3_2_constprop_o_ap_vld;

    assign l_TColl_2_3_3_constprop_o_ap_vld = grp_detectCollNode_fu_1055_l_TColl_2_3_3_constprop_o_ap_vld;

    assign numVertices_2_fu_1815_p2 = (numVertices_1_reg_2362 + 32'd1);

    assign or_ln110_fu_1610_p2 = (icmp_ln110_reg_2417 | icmp_ln110_1_reg_2422);

    assign or_ln119_fu_1761_p2 = (icmp_ln119_fu_1749_p2 | icmp_ln119_1_fu_1755_p2);

    assign or_ln138_fu_1956_p2 = (icmp_ln138_reg_2511 | icmp_ln138_1_reg_2516);

    assign or_ln188_fu_1803_p2 = (icmp_ln188_fu_1791_p2 | icmp_ln188_1_fu_1797_p2);

    assign p_shl1_fu_1867_p3 = {{select_ln96_5_reg_2492}, {3'd0}};

    assign p_shl_fu_1672_p3 = {{select_ln96_reg_2439}, {3'd0}};

    assign rand_int_fu_1564_p3 = {{xor_ln38_reg_2391}, {lshr_ln_reg_2386}};

    assign select_ln96_5_fu_1859_p3 = ((icmp35_fu_1847_p2[0:0] == 1'b1) ? add_ln96_fu_1853_p2 : 32'd0);

    assign select_ln96_fu_1664_p3 = ((icmp_fu_1653_p2[0:0] == 1'b1) ? add_ln96_2_fu_1659_p2 : 32'd0);

    assign sub_ln114_fu_1720_p2 = (tmp_26_fu_1704_p3 - tmp_27_fu_1712_p3);

    assign sub_ln130_fu_1634_p2 = (tmp_fu_1620_p3 - tmp_24_fu_1627_p3);

    assign sub_ln139_fu_1980_p2 = (tmp_35_fu_1966_p3 - tmp_36_fu_1973_p3);

    assign sub_ln294_fu_1915_p2 = (tmp_31_fu_1899_p3 - tmp_32_fu_1907_p3);

    assign sub_ln296_1_fu_1885_p2 = (p_shl1_fu_1867_p3 - zext_ln296_1_fu_1881_p1);

    assign sub_ln296_fu_1690_p2 = (p_shl_fu_1672_p3 - zext_ln296_fu_1686_p1);

    assign this_0_0_0_0_address0 = grp_detectCollNode_fu_1055_this_env_0_0_0_address0;

    assign this_0_0_0_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_0_0_ce0;

    assign this_0_0_0_1_address0 = grp_detectCollNode_fu_1055_this_env_0_0_1_address0;

    assign this_0_0_0_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_0_1_ce0;

    assign this_0_0_0_2_address0 = grp_detectCollNode_fu_1055_this_env_0_0_2_address0;

    assign this_0_0_0_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_0_2_ce0;

    assign this_0_0_1_0_address0 = grp_detectCollNode_fu_1055_this_env_0_1_0_address0;

    assign this_0_0_1_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_1_0_ce0;

    assign this_0_0_1_1_address0 = grp_detectCollNode_fu_1055_this_env_0_1_1_address0;

    assign this_0_0_1_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_1_1_ce0;

    assign this_0_0_1_2_address0 = grp_detectCollNode_fu_1055_this_env_0_1_2_address0;

    assign this_0_0_1_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_1_2_ce0;

    assign this_0_0_2_0_address0 = grp_detectCollNode_fu_1055_this_env_0_2_0_address0;

    assign this_0_0_2_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_2_0_ce0;

    assign this_0_0_2_1_address0 = grp_detectCollNode_fu_1055_this_env_0_2_1_address0;

    assign this_0_0_2_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_2_1_ce0;

    assign this_0_0_2_2_address0 = grp_detectCollNode_fu_1055_this_env_0_2_2_address0;

    assign this_0_0_2_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_2_2_ce0;

    assign this_0_0_3_0_address0 = grp_detectCollNode_fu_1055_this_env_0_3_0_address0;

    assign this_0_0_3_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_3_0_ce0;

    assign this_0_0_3_1_address0 = grp_detectCollNode_fu_1055_this_env_0_3_1_address0;

    assign this_0_0_3_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_3_1_ce0;

    assign this_0_0_3_2_address0 = grp_detectCollNode_fu_1055_this_env_0_3_2_address0;

    assign this_0_0_3_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_3_2_ce0;

    assign this_0_0_4_0_address0 = grp_detectCollNode_fu_1055_this_env_0_4_0_address0;

    assign this_0_0_4_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_4_0_ce0;

    assign this_0_0_4_1_address0 = grp_detectCollNode_fu_1055_this_env_0_4_1_address0;

    assign this_0_0_4_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_4_1_ce0;

    assign this_0_0_4_2_address0 = grp_detectCollNode_fu_1055_this_env_0_4_2_address0;

    assign this_0_0_4_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_4_2_ce0;

    assign this_0_0_5_0_address0 = grp_detectCollNode_fu_1055_this_env_0_5_0_address0;

    assign this_0_0_5_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_5_0_ce0;

    assign this_0_0_5_1_address0 = grp_detectCollNode_fu_1055_this_env_0_5_1_address0;

    assign this_0_0_5_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_5_1_ce0;

    assign this_0_0_5_2_address0 = grp_detectCollNode_fu_1055_this_env_0_5_2_address0;

    assign this_0_0_5_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_5_2_ce0;

    assign this_0_0_6_0_address0 = grp_detectCollNode_fu_1055_this_env_0_6_0_address0;

    assign this_0_0_6_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_6_0_ce0;

    assign this_0_0_6_1_address0 = grp_detectCollNode_fu_1055_this_env_0_6_1_address0;

    assign this_0_0_6_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_6_1_ce0;

    assign this_0_0_6_2_address0 = grp_detectCollNode_fu_1055_this_env_0_6_2_address0;

    assign this_0_0_6_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_6_2_ce0;

    assign this_0_0_7_0_address0 = grp_detectCollNode_fu_1055_this_env_0_7_0_address0;

    assign this_0_0_7_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_7_0_ce0;

    assign this_0_0_7_1_address0 = grp_detectCollNode_fu_1055_this_env_0_7_1_address0;

    assign this_0_0_7_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_7_1_ce0;

    assign this_0_0_7_2_address0 = grp_detectCollNode_fu_1055_this_env_0_7_2_address0;

    assign this_0_0_7_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_7_2_ce0;

    assign this_0_0_8_0_address0 = grp_detectCollNode_fu_1055_this_env_0_8_0_address0;

    assign this_0_0_8_0_ce0 = grp_detectCollNode_fu_1055_this_env_0_8_0_ce0;

    assign this_0_0_8_1_address0 = grp_detectCollNode_fu_1055_this_env_0_8_1_address0;

    assign this_0_0_8_1_ce0 = grp_detectCollNode_fu_1055_this_env_0_8_1_ce0;

    assign this_0_0_8_2_address0 = grp_detectCollNode_fu_1055_this_env_0_8_2_address0;

    assign this_0_0_8_2_ce0 = grp_detectCollNode_fu_1055_this_env_0_8_2_ce0;

    assign this_0_1_address0 = grp_detectCollNode_fu_1055_this_env_1_address0;

    assign this_0_1_address1 = grp_detectCollNode_fu_1055_this_env_1_address1;

    assign this_0_1_ce0 = grp_detectCollNode_fu_1055_this_env_1_ce0;

    assign this_0_1_ce1 = grp_detectCollNode_fu_1055_this_env_1_ce1;

    assign this_15_address0 = grp_detectCollNode_fu_1055_this_cPoints_address0;

    assign this_15_address1 = grp_detectCollNode_fu_1055_this_cPoints_address1;

    assign this_15_ce0 = grp_detectCollNode_fu_1055_this_cPoints_ce0;

    assign this_15_ce1 = grp_detectCollNode_fu_1055_this_cPoints_ce1;

    assign this_15_d0 = grp_detectCollNode_fu_1055_this_cPoints_d0;

    assign this_15_d1 = grp_detectCollNode_fu_1055_this_cPoints_d1;

    assign this_15_we0 = grp_detectCollNode_fu_1055_this_cPoints_we0;

    assign this_15_we1 = grp_detectCollNode_fu_1055_this_cPoints_we1;

    assign this_16_address0 = grp_detectCollNode_fu_1055_this_cAxes_address0;

    assign this_16_address1 = grp_detectCollNode_fu_1055_this_cAxes_address1;

    assign this_16_ce0 = grp_detectCollNode_fu_1055_this_cAxes_ce0;

    assign this_16_ce1 = grp_detectCollNode_fu_1055_this_cAxes_ce1;

    assign this_16_d0 = grp_detectCollNode_fu_1055_this_cAxes_d0;

    assign this_16_we0 = grp_detectCollNode_fu_1055_this_cAxes_we0;

    assign this_4_0_0_address0 = grp_detectCollNode_fu_1055_this_TLink_0_0_address0;

    assign this_4_0_0_ce0 = grp_detectCollNode_fu_1055_this_TLink_0_0_ce0;

    assign this_4_0_1_address0 = grp_detectCollNode_fu_1055_this_TLink_0_1_address0;

    assign this_4_0_1_ce0 = grp_detectCollNode_fu_1055_this_TLink_0_1_ce0;

    assign this_4_0_2_address0 = grp_detectCollNode_fu_1055_this_TLink_0_2_address0;

    assign this_4_0_2_ce0 = grp_detectCollNode_fu_1055_this_TLink_0_2_ce0;

    assign this_4_0_3_address0 = grp_detectCollNode_fu_1055_this_TLink_0_3_address0;

    assign this_4_0_3_ce0 = grp_detectCollNode_fu_1055_this_TLink_0_3_ce0;

    assign this_4_1_0_address0 = grp_detectCollNode_fu_1055_this_TLink_1_0_address0;

    assign this_4_1_0_ce0 = grp_detectCollNode_fu_1055_this_TLink_1_0_ce0;

    assign this_4_1_1_address0 = grp_detectCollNode_fu_1055_this_TLink_1_1_address0;

    assign this_4_1_1_ce0 = grp_detectCollNode_fu_1055_this_TLink_1_1_ce0;

    assign this_4_1_2_address0 = grp_detectCollNode_fu_1055_this_TLink_1_2_address0;

    assign this_4_1_2_ce0 = grp_detectCollNode_fu_1055_this_TLink_1_2_ce0;

    assign this_4_1_3_address0 = grp_detectCollNode_fu_1055_this_TLink_1_3_address0;

    assign this_4_1_3_ce0 = grp_detectCollNode_fu_1055_this_TLink_1_3_ce0;

    assign this_4_2_0_address0 = grp_detectCollNode_fu_1055_this_TLink_2_0_address0;

    assign this_4_2_0_ce0 = grp_detectCollNode_fu_1055_this_TLink_2_0_ce0;

    assign this_4_2_1_address0 = grp_detectCollNode_fu_1055_this_TLink_2_1_address0;

    assign this_4_2_1_ce0 = grp_detectCollNode_fu_1055_this_TLink_2_1_ce0;

    assign this_4_2_2_address0 = grp_detectCollNode_fu_1055_this_TLink_2_2_address0;

    assign this_4_2_2_ce0 = grp_detectCollNode_fu_1055_this_TLink_2_2_ce0;

    assign this_4_2_3_address0 = grp_detectCollNode_fu_1055_this_TLink_2_3_address0;

    assign this_4_2_3_ce0 = grp_detectCollNode_fu_1055_this_TLink_2_3_ce0;

    assign this_4_3_0_address0 = grp_detectCollNode_fu_1055_this_TLink_3_0_address0;

    assign this_4_3_0_ce0 = grp_detectCollNode_fu_1055_this_TLink_3_0_ce0;

    assign this_4_3_1_address0 = grp_detectCollNode_fu_1055_this_TLink_3_1_address0;

    assign this_4_3_1_ce0 = grp_detectCollNode_fu_1055_this_TLink_3_1_ce0;

    assign this_4_3_2_address0 = grp_detectCollNode_fu_1055_this_TLink_3_2_address0;

    assign this_4_3_2_ce0 = grp_detectCollNode_fu_1055_this_TLink_3_2_ce0;

    assign this_4_3_3_address0 = grp_detectCollNode_fu_1055_this_TLink_3_3_address0;

    assign this_4_3_3_ce0 = grp_detectCollNode_fu_1055_this_TLink_3_3_ce0;

    assign this_5_0_0_address0 = grp_detectCollNode_fu_1055_this_TJoint_0_0_address0;

    assign this_5_0_0_ce0 = grp_detectCollNode_fu_1055_this_TJoint_0_0_ce0;

    assign this_5_0_0_d0 = grp_detectCollNode_fu_1055_this_TJoint_0_0_d0;

    assign this_5_0_0_we0 = grp_detectCollNode_fu_1055_this_TJoint_0_0_we0;

    assign this_5_0_1_address0 = grp_detectCollNode_fu_1055_this_TJoint_0_1_address0;

    assign this_5_0_1_ce0 = grp_detectCollNode_fu_1055_this_TJoint_0_1_ce0;

    assign this_5_0_1_d0 = grp_detectCollNode_fu_1055_this_TJoint_0_1_d0;

    assign this_5_0_1_we0 = grp_detectCollNode_fu_1055_this_TJoint_0_1_we0;

    assign this_5_0_2_address0 = grp_detectCollNode_fu_1055_this_TJoint_0_2_address0;

    assign this_5_0_2_ce0 = grp_detectCollNode_fu_1055_this_TJoint_0_2_ce0;

    assign this_5_0_2_d0 = grp_detectCollNode_fu_1055_this_TJoint_0_2_d0;

    assign this_5_0_2_we0 = grp_detectCollNode_fu_1055_this_TJoint_0_2_we0;

    assign this_5_0_3_address0 = grp_detectCollNode_fu_1055_this_TJoint_0_3_address0;

    assign this_5_0_3_ce0 = grp_detectCollNode_fu_1055_this_TJoint_0_3_ce0;

    assign this_5_0_3_d0 = grp_detectCollNode_fu_1055_this_TJoint_0_3_d0;

    assign this_5_0_3_we0 = grp_detectCollNode_fu_1055_this_TJoint_0_3_we0;

    assign this_5_1_0_address0 = grp_detectCollNode_fu_1055_this_TJoint_1_0_address0;

    assign this_5_1_0_ce0 = grp_detectCollNode_fu_1055_this_TJoint_1_0_ce0;

    assign this_5_1_0_d0 = grp_detectCollNode_fu_1055_this_TJoint_1_0_d0;

    assign this_5_1_0_we0 = grp_detectCollNode_fu_1055_this_TJoint_1_0_we0;

    assign this_5_1_1_address0 = grp_detectCollNode_fu_1055_this_TJoint_1_1_address0;

    assign this_5_1_1_ce0 = grp_detectCollNode_fu_1055_this_TJoint_1_1_ce0;

    assign this_5_1_1_d0 = grp_detectCollNode_fu_1055_this_TJoint_1_1_d0;

    assign this_5_1_1_we0 = grp_detectCollNode_fu_1055_this_TJoint_1_1_we0;

    assign this_5_1_2_address0 = grp_detectCollNode_fu_1055_this_TJoint_1_2_address0;

    assign this_5_1_2_ce0 = grp_detectCollNode_fu_1055_this_TJoint_1_2_ce0;

    assign this_5_1_2_d0 = grp_detectCollNode_fu_1055_this_TJoint_1_2_d0;

    assign this_5_1_2_we0 = grp_detectCollNode_fu_1055_this_TJoint_1_2_we0;

    assign this_5_1_3_address0 = grp_detectCollNode_fu_1055_this_TJoint_1_3_address0;

    assign this_5_1_3_ce0 = grp_detectCollNode_fu_1055_this_TJoint_1_3_ce0;

    assign this_5_1_3_d0 = grp_detectCollNode_fu_1055_this_TJoint_1_3_d0;

    assign this_5_1_3_we0 = grp_detectCollNode_fu_1055_this_TJoint_1_3_we0;

    assign this_5_2_0_address0 = grp_detectCollNode_fu_1055_this_TJoint_2_0_address0;

    assign this_5_2_0_ce0 = grp_detectCollNode_fu_1055_this_TJoint_2_0_ce0;

    assign this_5_2_0_d0 = grp_detectCollNode_fu_1055_this_TJoint_2_0_d0;

    assign this_5_2_0_we0 = grp_detectCollNode_fu_1055_this_TJoint_2_0_we0;

    assign this_5_2_1_address0 = grp_detectCollNode_fu_1055_this_TJoint_2_1_address0;

    assign this_5_2_1_ce0 = grp_detectCollNode_fu_1055_this_TJoint_2_1_ce0;

    assign this_5_2_1_d0 = grp_detectCollNode_fu_1055_this_TJoint_2_1_d0;

    assign this_5_2_1_we0 = grp_detectCollNode_fu_1055_this_TJoint_2_1_we0;

    assign this_5_2_2_address0 = grp_detectCollNode_fu_1055_this_TJoint_2_2_address0;

    assign this_5_2_2_ce0 = grp_detectCollNode_fu_1055_this_TJoint_2_2_ce0;

    assign this_5_2_2_d0 = grp_detectCollNode_fu_1055_this_TJoint_2_2_d0;

    assign this_5_2_2_we0 = grp_detectCollNode_fu_1055_this_TJoint_2_2_we0;

    assign this_5_2_3_address0 = grp_detectCollNode_fu_1055_this_TJoint_2_3_address0;

    assign this_5_2_3_ce0 = grp_detectCollNode_fu_1055_this_TJoint_2_3_ce0;

    assign this_5_2_3_d0 = grp_detectCollNode_fu_1055_this_TJoint_2_3_d0;

    assign this_5_2_3_we0 = grp_detectCollNode_fu_1055_this_TJoint_2_3_we0;

    assign this_5_3_0_address0 = grp_detectCollNode_fu_1055_this_TJoint_3_0_address0;

    assign this_5_3_0_ce0 = grp_detectCollNode_fu_1055_this_TJoint_3_0_ce0;

    assign this_5_3_0_d0 = grp_detectCollNode_fu_1055_this_TJoint_3_0_d0;

    assign this_5_3_0_we0 = grp_detectCollNode_fu_1055_this_TJoint_3_0_we0;

    assign this_5_3_1_address0 = grp_detectCollNode_fu_1055_this_TJoint_3_1_address0;

    assign this_5_3_1_ce0 = grp_detectCollNode_fu_1055_this_TJoint_3_1_ce0;

    assign this_5_3_1_d0 = grp_detectCollNode_fu_1055_this_TJoint_3_1_d0;

    assign this_5_3_1_we0 = grp_detectCollNode_fu_1055_this_TJoint_3_1_we0;

    assign this_5_3_2_address0 = grp_detectCollNode_fu_1055_this_TJoint_3_2_address0;

    assign this_5_3_2_ce0 = grp_detectCollNode_fu_1055_this_TJoint_3_2_ce0;

    assign this_5_3_2_d0 = grp_detectCollNode_fu_1055_this_TJoint_3_2_d0;

    assign this_5_3_2_we0 = grp_detectCollNode_fu_1055_this_TJoint_3_2_we0;

    assign this_5_3_3_address0 = grp_detectCollNode_fu_1055_this_TJoint_3_3_address0;

    assign this_5_3_3_ce0 = grp_detectCollNode_fu_1055_this_TJoint_3_3_ce0;

    assign this_5_3_3_d0 = grp_detectCollNode_fu_1055_this_TJoint_3_3_d0;

    assign this_5_3_3_we0 = grp_detectCollNode_fu_1055_this_TJoint_3_3_we0;

    assign this_6_0_0_address0 = grp_detectCollNode_fu_1055_this_TCurr_0_0_address0;

    assign this_6_0_0_ce0 = grp_detectCollNode_fu_1055_this_TCurr_0_0_ce0;

    assign this_6_0_0_d0 = grp_detectCollNode_fu_1055_this_TCurr_0_0_d0;

    assign this_6_0_0_we0 = grp_detectCollNode_fu_1055_this_TCurr_0_0_we0;

    assign this_6_0_1_address0 = grp_detectCollNode_fu_1055_this_TCurr_0_1_address0;

    assign this_6_0_1_ce0 = grp_detectCollNode_fu_1055_this_TCurr_0_1_ce0;

    assign this_6_0_1_d0 = grp_detectCollNode_fu_1055_this_TCurr_0_1_d0;

    assign this_6_0_1_we0 = grp_detectCollNode_fu_1055_this_TCurr_0_1_we0;

    assign this_6_0_2_address0 = grp_detectCollNode_fu_1055_this_TCurr_0_2_address0;

    assign this_6_0_2_ce0 = grp_detectCollNode_fu_1055_this_TCurr_0_2_ce0;

    assign this_6_0_2_d0 = grp_detectCollNode_fu_1055_this_TCurr_0_2_d0;

    assign this_6_0_2_we0 = grp_detectCollNode_fu_1055_this_TCurr_0_2_we0;

    assign this_6_0_3_address0 = grp_detectCollNode_fu_1055_this_TCurr_0_3_address0;

    assign this_6_0_3_ce0 = grp_detectCollNode_fu_1055_this_TCurr_0_3_ce0;

    assign this_6_0_3_d0 = grp_detectCollNode_fu_1055_this_TCurr_0_3_d0;

    assign this_6_0_3_we0 = grp_detectCollNode_fu_1055_this_TCurr_0_3_we0;

    assign this_6_1_0_address0 = grp_detectCollNode_fu_1055_this_TCurr_1_0_address0;

    assign this_6_1_0_ce0 = grp_detectCollNode_fu_1055_this_TCurr_1_0_ce0;

    assign this_6_1_0_d0 = grp_detectCollNode_fu_1055_this_TCurr_1_0_d0;

    assign this_6_1_0_we0 = grp_detectCollNode_fu_1055_this_TCurr_1_0_we0;

    assign this_6_1_1_address0 = grp_detectCollNode_fu_1055_this_TCurr_1_1_address0;

    assign this_6_1_1_ce0 = grp_detectCollNode_fu_1055_this_TCurr_1_1_ce0;

    assign this_6_1_1_d0 = grp_detectCollNode_fu_1055_this_TCurr_1_1_d0;

    assign this_6_1_1_we0 = grp_detectCollNode_fu_1055_this_TCurr_1_1_we0;

    assign this_6_1_2_address0 = grp_detectCollNode_fu_1055_this_TCurr_1_2_address0;

    assign this_6_1_2_ce0 = grp_detectCollNode_fu_1055_this_TCurr_1_2_ce0;

    assign this_6_1_2_d0 = grp_detectCollNode_fu_1055_this_TCurr_1_2_d0;

    assign this_6_1_2_we0 = grp_detectCollNode_fu_1055_this_TCurr_1_2_we0;

    assign this_6_1_3_address0 = grp_detectCollNode_fu_1055_this_TCurr_1_3_address0;

    assign this_6_1_3_ce0 = grp_detectCollNode_fu_1055_this_TCurr_1_3_ce0;

    assign this_6_1_3_d0 = grp_detectCollNode_fu_1055_this_TCurr_1_3_d0;

    assign this_6_1_3_we0 = grp_detectCollNode_fu_1055_this_TCurr_1_3_we0;

    assign this_6_2_0_address0 = grp_detectCollNode_fu_1055_this_TCurr_2_0_address0;

    assign this_6_2_0_ce0 = grp_detectCollNode_fu_1055_this_TCurr_2_0_ce0;

    assign this_6_2_0_d0 = grp_detectCollNode_fu_1055_this_TCurr_2_0_d0;

    assign this_6_2_0_we0 = grp_detectCollNode_fu_1055_this_TCurr_2_0_we0;

    assign this_6_2_1_address0 = grp_detectCollNode_fu_1055_this_TCurr_2_1_address0;

    assign this_6_2_1_ce0 = grp_detectCollNode_fu_1055_this_TCurr_2_1_ce0;

    assign this_6_2_1_d0 = grp_detectCollNode_fu_1055_this_TCurr_2_1_d0;

    assign this_6_2_1_we0 = grp_detectCollNode_fu_1055_this_TCurr_2_1_we0;

    assign this_6_2_2_address0 = grp_detectCollNode_fu_1055_this_TCurr_2_2_address0;

    assign this_6_2_2_ce0 = grp_detectCollNode_fu_1055_this_TCurr_2_2_ce0;

    assign this_6_2_2_d0 = grp_detectCollNode_fu_1055_this_TCurr_2_2_d0;

    assign this_6_2_2_we0 = grp_detectCollNode_fu_1055_this_TCurr_2_2_we0;

    assign this_6_2_3_address0 = grp_detectCollNode_fu_1055_this_TCurr_2_3_address0;

    assign this_6_2_3_ce0 = grp_detectCollNode_fu_1055_this_TCurr_2_3_ce0;

    assign this_6_2_3_d0 = grp_detectCollNode_fu_1055_this_TCurr_2_3_d0;

    assign this_6_2_3_we0 = grp_detectCollNode_fu_1055_this_TCurr_2_3_we0;

    assign this_6_3_0_address0 = grp_detectCollNode_fu_1055_this_TCurr_3_0_address0;

    assign this_6_3_0_ce0 = grp_detectCollNode_fu_1055_this_TCurr_3_0_ce0;

    assign this_6_3_0_d0 = grp_detectCollNode_fu_1055_this_TCurr_3_0_d0;

    assign this_6_3_0_we0 = grp_detectCollNode_fu_1055_this_TCurr_3_0_we0;

    assign this_6_3_1_address0 = grp_detectCollNode_fu_1055_this_TCurr_3_1_address0;

    assign this_6_3_1_ce0 = grp_detectCollNode_fu_1055_this_TCurr_3_1_ce0;

    assign this_6_3_1_d0 = grp_detectCollNode_fu_1055_this_TCurr_3_1_d0;

    assign this_6_3_1_we0 = grp_detectCollNode_fu_1055_this_TCurr_3_1_we0;

    assign this_6_3_2_address0 = grp_detectCollNode_fu_1055_this_TCurr_3_2_address0;

    assign this_6_3_2_ce0 = grp_detectCollNode_fu_1055_this_TCurr_3_2_ce0;

    assign this_6_3_2_d0 = grp_detectCollNode_fu_1055_this_TCurr_3_2_d0;

    assign this_6_3_2_we0 = grp_detectCollNode_fu_1055_this_TCurr_3_2_we0;

    assign this_6_3_3_address0 = grp_detectCollNode_fu_1055_this_TCurr_3_3_address0;

    assign this_6_3_3_ce0 = grp_detectCollNode_fu_1055_this_TCurr_3_3_ce0;

    assign this_6_3_3_d0 = grp_detectCollNode_fu_1055_this_TCurr_3_3_d0;

    assign this_6_3_3_we0 = grp_detectCollNode_fu_1055_this_TCurr_3_3_we0;

    assign this_7_address0 = grp_detectCollNode_fu_1055_this_q_address0;

    assign this_7_ce0 = grp_detectCollNode_fu_1055_this_q_ce0;

    assign this_7_d0 = grp_detectCollNode_fu_1055_this_q_d0;

    assign this_7_we0 = grp_detectCollNode_fu_1055_this_q_we0;

    assign tmp_16_fu_1512_p3 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out[32'd3];

    assign tmp_17_fu_1520_p3 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out[32'd5];

    assign tmp_18_fu_1528_p3 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_or_i_i_i110_out[32'd2];

    assign tmp_19_fu_1644_p4 = {{numVertices_1_reg_2362[31:1]}};

    assign tmp_20_fu_1837_p4 = {{numVertices_fu_520[31:1]}};

    assign tmp_24_fu_1627_p3 = {{trunc_ln83_reg_2369}, {1'd0}};

    assign tmp_25_fu_1679_p3 = {{select_ln96_reg_2439}, {1'd0}};

    assign tmp_262_fu_1584_p4 = {{bitcast_ln110_fu_1581_p1[62:52]}};

    assign tmp_264_fu_1735_p4 = {{bitcast_ln119_fu_1731_p1[62:52]}};

    assign tmp_266_fu_1777_p4 = {{bitcast_ln188_fu_1773_p1[62:52]}};

    assign tmp_268_fu_1930_p4 = {{bitcast_ln138_fu_1926_p1[62:52]}};

    assign tmp_26_fu_1704_p3 = {{empty_fu_1700_p1}, {3'd0}};

    assign tmp_27_fu_1712_p3 = {{bestIdx_3_loc_fu_540}, {1'd0}};

    assign tmp_30_fu_1874_p3 = {{select_ln96_5_reg_2492}, {1'd0}};

    assign tmp_31_fu_1899_p3 = {{empty_64_fu_1895_p1}, {3'd0}};

    assign tmp_32_fu_1907_p3 = {{bestIdx_6_loc_fu_528}, {1'd0}};

    assign tmp_35_fu_1966_p3 = {{trunc_ln83_3_reg_2487}, {3'd0}};

    assign tmp_36_fu_1973_p3 = {{trunc_ln83_2_reg_2482}, {1'd0}};

    assign tmp_fu_1620_p3 = {{trunc_ln83_1_reg_2374}, {3'd0}};

    assign trunc_ln110_fu_1594_p1 = bitcast_ln110_fu_1581_p1[51:0];

    assign trunc_ln119_fu_1745_p1 = bitcast_ln119_fu_1731_p1[51:0];

    assign trunc_ln138_fu_1940_p1 = bitcast_ln138_fu_1926_p1[51:0];

    assign trunc_ln188_fu_1787_p1 = bitcast_ln188_fu_1773_p1[51:0];

    assign trunc_ln37_fu_1508_p1 = grp_planRRT_Pipeline_VITIS_LOOP_152_1_fu_980_shr6_i_i_i_phi_out[0:0];

    assign trunc_ln83_1_fu_1487_p1 = numVertices_fu_520[9:0];

    assign trunc_ln83_2_fu_1829_p1 = numVertices_fu_520[11:0];

    assign trunc_ln83_3_fu_1833_p1 = numVertices_fu_520[9:0];

    assign trunc_ln83_fu_1483_p1 = numVertices_fu_520[11:0];

    assign xor_ln38_2_fu_1546_p2 = (trunc_ln37_fu_1508_p1 ^ tmp_16_fu_1512_p3);

    assign xor_ln38_3_fu_1552_p2 = (tmp_18_fu_1528_p3 ^ tmp_17_fu_1520_p3);

    assign xor_ln38_fu_1558_p2 = (xor_ln38_3_fu_1552_p2 ^ xor_ln38_2_fu_1546_p2);

    assign zext_ln296_1_fu_1881_p1 = tmp_30_fu_1874_p3;

    assign zext_ln296_fu_1686_p1 = tmp_25_fu_1679_p3;

    assign zext_ln47_fu_1576_p1 = rand_int_fu_1564_p3;

    always @(posedge ap_clk) begin
        sub_ln130_reg_2431[0]   <= 1'b0;
        sub_ln296_reg_2445[0]   <= 1'b0;
        sub_ln114_reg_2450[0]   <= 1'b0;
        sub_ln296_1_reg_2498[0] <= 1'b0;
        sub_ln294_reg_2503[0]   <= 1'b0;
        sub_ln139_reg_2524[0]   <= 1'b0;
    end

endmodule  //main_planRRT
