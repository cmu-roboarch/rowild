/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_atan2_generic_double_Pipeline_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    y_1,
    zext_ln681,
    z_out,
    z_out_ap_vld
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [88:0] y_1;
    input [85:0] zext_ln681;
    output [85:0] z_out;
    output z_out_ap_vld;

    reg ap_idle;
    reg z_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln138_fu_139_p2;
    reg    ap_condition_exit_pp0_iter1_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire   [6:0] cordic_ctab_table_128_address0;
    reg    cordic_ctab_table_128_ce0;
    wire   [125:0] cordic_ctab_table_128_q0;
    wire    ap_block_pp0_stage0_11001;
    reg   [0:0] icmp_ln138_reg_331;
    wire   [0:0] tmp_fu_162_p3;
    reg   [0:0] tmp_reg_335;
    reg   [0:0] tmp_reg_335_pp0_iter2_reg;
    reg   [84:0] trunc_ln_reg_345;
    reg   [0:0] tmp_27_reg_350;
    wire   [63:0] zext_ln138_fu_157_p1;
    wire    ap_block_pp0_stage0;
    reg   [88:0] x_fu_64;
    wire   [88:0] x_2_fu_192_p3;
    wire   [88:0] zext_ln681_cast_fu_112_p1;
    wire    ap_loop_init;
    reg   [88:0] y_fu_68;
    wire   [88:0] y_2_fu_218_p3;
    reg   [85:0] z_fu_72;
    wire   [85:0] z_1_fu_286_p3;
    reg   [6:0] k_fu_76;
    wire   [6:0] add_ln138_fu_145_p2;
    wire    ap_block_pp0_stage0_01001;
    wire   [88:0] zext_ln159_fu_170_p1;
    wire   [88:0] y_s_fu_174_p2;
    wire   [88:0] sub_ln101_fu_180_p2;
    wire   [88:0] add_ln101_fu_186_p2;
    wire   [88:0] x_s_fu_200_p2;
    wire   [88:0] add_ln101_1_fu_212_p2;
    wire   [88:0] sub_ln101_1_fu_206_p2;
    wire   [84:0] zext_ln163_fu_262_p1;
    wire   [84:0] add_ln163_fu_265_p2;
    wire   [85:0] zext_ln164_fu_270_p1;
    wire   [85:0] sub_ln101_2_fu_274_p2;
    wire   [85:0] add_ln101_2_fu_280_p2;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 x_fu_64 = 89'd0;
        #0 y_fu_68 = 89'd0;
        #0 z_fu_72 = 86'd0;
        #0 k_fu_76 = 7'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_atan2_generic_double_Pipeline_1_cordic_ctab_table_128_ROM_AUTO_1R #(
        .DataWidth(126),
        .AddressRange(128),
        .AddressWidth(7)
    ) cordic_ctab_table_128_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(cordic_ctab_table_128_address0),
        .ce0(cordic_ctab_table_128_ce0),
        .q0(cordic_ctab_table_128_q0)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
                ap_enable_reg_pp0_iter2 <= 1'b0;
            end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                k_fu_76 <= 7'd0;
            end else if (((icmp_ln138_fu_139_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                k_fu_76 <= add_ln138_fu_145_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                x_fu_64 <= zext_ln681_cast_fu_112_p1;
            end else if (((icmp_ln138_fu_139_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                x_fu_64 <= x_2_fu_192_p3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                y_fu_68 <= y_1;
            end else if (((icmp_ln138_fu_139_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                y_fu_68 <= y_2_fu_218_p3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                z_fu_72 <= 86'd0;
            end else if ((ap_enable_reg_pp0_iter3 == 1'b1)) begin
                z_fu_72 <= z_1_fu_286_p3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
            icmp_ln138_reg_331 <= icmp_ln138_fu_139_p2;
            tmp_reg_335 <= y_fu_68[32'd88];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            tmp_27_reg_350 <= cordic_ctab_table_128_q0[32'd40];
            tmp_reg_335_pp0_iter2_reg <= tmp_reg_335;
            trunc_ln_reg_345 <= {{cordic_ctab_table_128_q0[125:41]}};
        end
    end

    always @(*) begin
        if (((icmp_ln138_fu_139_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter1_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter1_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            cordic_ctab_table_128_ce0 = 1'b1;
        end else begin
            cordic_ctab_table_128_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln138_reg_331 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            z_out_ap_vld = 1'b1;
        end else begin
            z_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln101_1_fu_212_p2 = (x_s_fu_200_p2 + y_fu_68);

    assign add_ln101_2_fu_280_p2 = (zext_ln164_fu_270_p1 + z_fu_72);

    assign add_ln101_fu_186_p2 = (y_s_fu_174_p2 + x_fu_64);

    assign add_ln138_fu_145_p2 = (k_fu_76 + 7'd1);

    assign add_ln163_fu_265_p2 = (zext_ln163_fu_262_p1 + trunc_ln_reg_345);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

    assign cordic_ctab_table_128_address0 = zext_ln138_fu_157_p1;

    assign icmp_ln138_fu_139_p2 = ((k_fu_76 == 7'd88) ? 1'b1 : 1'b0);

    assign sub_ln101_1_fu_206_p2 = (y_fu_68 - x_s_fu_200_p2);

    assign sub_ln101_2_fu_274_p2 = (z_fu_72 - zext_ln164_fu_270_p1);

    assign sub_ln101_fu_180_p2 = (x_fu_64 - y_s_fu_174_p2);

    assign tmp_fu_162_p3 = y_fu_68[32'd88];

    assign x_2_fu_192_p3 = ((tmp_fu_162_p3[0:0] == 1'b1) ? sub_ln101_fu_180_p2 : add_ln101_fu_186_p2);

    assign x_s_fu_200_p2 = $signed(x_fu_64) >>> zext_ln159_fu_170_p1;

    assign y_2_fu_218_p3 = ((tmp_fu_162_p3[0:0] == 1'b1) ? add_ln101_1_fu_212_p2 : sub_ln101_1_fu_206_p2);

    assign y_s_fu_174_p2 = $signed(y_fu_68) >>> zext_ln159_fu_170_p1;

    assign z_1_fu_286_p3 = ((tmp_reg_335_pp0_iter2_reg[0:0] == 1'b1) ? sub_ln101_2_fu_274_p2 : add_ln101_2_fu_280_p2);

    assign z_out = z_fu_72;

    assign zext_ln138_fu_157_p1 = k_fu_76;

    assign zext_ln159_fu_170_p1 = k_fu_76;

    assign zext_ln163_fu_262_p1 = tmp_27_reg_350;

    assign zext_ln164_fu_270_p1 = add_ln163_fu_265_p2;

    assign zext_ln681_cast_fu_112_p1 = zext_ln681;

endmodule  //main_atan2_generic_double_Pipeline_1
