/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    minDist_4,
    sub_ln296_1,
    rrtVertices_address0,
    rrtVertices_ce0,
    rrtVertices_q0,
    bestIdx_6_out,
    bestIdx_6_out_ap_vld,
    goal_address0,
    goal_ce0,
    goal_q0,
    grp_fu_2529_p_din0,
    grp_fu_2529_p_din1,
    grp_fu_2529_p_opcode,
    grp_fu_2529_p_dout0,
    grp_fu_2529_p_ce,
    grp_fu_2533_p_din0,
    grp_fu_2533_p_din1,
    grp_fu_2533_p_dout0,
    grp_fu_2533_p_ce,
    grp_fu_1454_p_din0,
    grp_fu_1454_p_din1,
    grp_fu_1454_p_opcode,
    grp_fu_1454_p_dout0,
    grp_fu_1454_p_ce,
    grp_fu_1462_p_din0,
    grp_fu_1462_p_din1,
    grp_fu_1462_p_dout0,
    grp_fu_1462_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 8'd1;
    parameter ap_ST_fsm_pp0_stage1 = 8'd2;
    parameter ap_ST_fsm_pp0_stage2 = 8'd4;
    parameter ap_ST_fsm_pp0_stage3 = 8'd8;
    parameter ap_ST_fsm_pp0_stage4 = 8'd16;
    parameter ap_ST_fsm_pp0_stage5 = 8'd32;
    parameter ap_ST_fsm_pp0_stage6 = 8'd64;
    parameter ap_ST_fsm_pp0_stage7 = 8'd128;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] minDist_4;
    input [34:0] sub_ln296_1;
    output [12:0] rrtVertices_address0;
    output rrtVertices_ce0;
    input [63:0] rrtVertices_q0;
    output [11:0] bestIdx_6_out;
    output bestIdx_6_out_ap_vld;
    output [2:0] goal_address0;
    output goal_ce0;
    input [63:0] goal_q0;
    output [63:0] grp_fu_2529_p_din0;
    output [63:0] grp_fu_2529_p_din1;
    output [1:0] grp_fu_2529_p_opcode;
    input [63:0] grp_fu_2529_p_dout0;
    output grp_fu_2529_p_ce;
    output [63:0] grp_fu_2533_p_din0;
    output [63:0] grp_fu_2533_p_din1;
    input [63:0] grp_fu_2533_p_dout0;
    output grp_fu_2533_p_ce;
    output [63:0] grp_fu_1454_p_din0;
    output [63:0] grp_fu_1454_p_din1;
    output [4:0] grp_fu_1454_p_opcode;
    input [0:0] grp_fu_1454_p_dout0;
    output grp_fu_1454_p_ce;
    output [63:0] grp_fu_1462_p_din0;
    output [63:0] grp_fu_1462_p_din1;
    input [63:0] grp_fu_1462_p_dout0;
    output grp_fu_1462_p_ce;

    reg ap_idle;
    reg rrtVertices_ce0;
    reg bestIdx_6_out_ap_vld;
    reg goal_ce0;

    (* fsm_encoding = "none" *) reg   [7:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_subdone;
    reg   [0:0] icmp_ln96_reg_499;
    reg    ap_condition_exit_pp0_iter0_stage7;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    reg   [30:0] idx_2_reg_489;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    reg   [30:0] idx_2_reg_489_pp0_iter1_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter2_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter3_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter4_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter5_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter6_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter7_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter8_reg;
    reg   [30:0] idx_2_reg_489_pp0_iter9_reg;
    reg   [34:0] indvar_flatten12_load_reg_494;
    wire   [0:0] icmp_ln96_fu_186_p2;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter1_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter2_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter3_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter4_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter5_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter6_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter7_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter8_reg;
    reg   [0:0] icmp_ln96_reg_499_pp0_iter9_reg;
    wire   [0:0] icmp_ln293_fu_200_p2;
    reg   [0:0] icmp_ln293_reg_503;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter1_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter2_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter3_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter4_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter5_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter6_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter7_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter8_reg;
    reg   [0:0] icmp_ln293_reg_503_pp0_iter9_reg;
    wire   [2:0] select_ln96_fu_206_p3;
    reg   [2:0] select_ln96_reg_510;
    wire   [12:0] add_ln294_fu_261_p2;
    reg   [12:0] add_ln294_reg_515;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [63:0] goal_load_reg_530;
    reg   [63:0] rrtVertices_load_reg_535;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    reg   [63:0] sub_i9_i1_reg_540;
    wire   [63:0] select_ln96_1_fu_300_p3;
    reg   [63:0] select_ln96_1_reg_551;
    reg   [63:0] mul_i10_i1_reg_556;
    reg   [63:0] dist_2_reg_561;
    reg   [63:0] d_reg_566;
    reg   [63:0] minDist_1_reg_573;
    reg   [31:0] bestIdx_1_reg_581;
    wire   [0:0] and_ln98_1_fu_397_p2;
    reg   [0:0] and_ln98_1_reg_586;
    wire   [31:0] bestIdx_3_fu_403_p3;
    reg   [31:0] bestIdx_3_reg_591;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage3_subdone;
    reg    ap_condition_exit_pp0_iter9_stage3;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_subdone;
    wire   [63:0] zext_ln293_fu_252_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln294_1_fu_272_p1;
    wire    ap_block_pp0_stage2;
    reg   [63:0] dist_fu_64;
    reg   [63:0] ap_sig_allocacmp_dist_1;
    wire    ap_loop_init;
    reg   [2:0] i_fu_68;
    wire   [2:0] add_ln293_fu_281_p2;
    reg   [31:0] bestIdx_fu_72;
    wire   [31:0] select_ln96_4_fu_427_p3;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_block_pp0_stage3;
    reg   [63:0] minDist_fu_76;
    wire   [63:0] select_ln96_3_fu_421_p3;
    reg   [30:0] idx_fu_80;
    wire   [30:0] select_ln96_2_fu_214_p3;
    reg   [34:0] indvar_flatten12_fu_84;
    wire   [34:0] add_ln96_fu_276_p2;
    wire    ap_block_pp0_stage3_01001;
    wire    ap_block_pp0_stage0;
    reg   [63:0] grp_fu_133_p0;
    reg   [63:0] grp_fu_133_p1;
    wire    ap_block_pp0_stage4;
    wire   [30:0] add_ln96_1_fu_194_p2;
    wire   [9:0] trunc_ln294_1_fu_226_p1;
    wire   [11:0] trunc_ln294_fu_222_p1;
    wire   [12:0] tmp_33_fu_230_p3;
    wire   [12:0] tmp_34_fu_238_p3;
    wire   [12:0] sub_ln294_fu_246_p2;
    wire   [12:0] zext_ln294_fu_257_p1;
    wire   [63:0] bitcast_ln98_fu_321_p1;
    wire   [63:0] bitcast_ln98_1_fu_338_p1;
    wire   [10:0] tmp_368_dup_fu_324_p4;
    wire   [51:0] trunc_ln98_fu_334_p1;
    wire   [0:0] icmp_ln98_1_fu_361_p2;
    wire   [0:0] icmp_ln98_fu_355_p2;
    wire   [10:0] tmp_369_dup_fu_341_p4;
    wire   [51:0] trunc_ln98_1_fu_351_p1;
    wire   [0:0] icmp_ln98_3_fu_379_p2;
    wire   [0:0] icmp_ln98_2_fu_373_p2;
    wire   [0:0] or_ln98_fu_367_p2;
    wire   [0:0] or_ln98_1_fu_385_p2;
    wire   [0:0] and_ln98_fu_391_p2;
    wire   [31:0] zext_ln96_fu_318_p1;
    wire   [63:0] minDist_6_fu_416_p3;
    reg   [1:0] grp_fu_133_opcode;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage4_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    wire    ap_block_pp0_stage7_11001;
    reg    ap_idle_pp0_0to8;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg   [7:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to9;
    reg    ap_done_pending_pp0;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 8'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 dist_fu_64 = 64'd0;
        #0 i_fu_68 = 3'd0;
        #0 bestIdx_fu_72 = 32'd0;
        #0 minDist_fu_76 = 64'd0;
        #0 idx_fu_80 = 31'd0;
        #0 indvar_flatten12_fu_84 = 35'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage7),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b1 == ap_condition_exit_pp0_iter9_stage3) | ((1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
                ap_enable_reg_pp0_iter9 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3)) | ((1'b0 == ap_block_pp0_stage4_subdone) & (ap_loop_exit_ready_pp0_iter8_reg == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            bestIdx_fu_72 <= 32'd0;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln96_reg_499_pp0_iter9_reg == 1'd0))) begin
            bestIdx_fu_72 <= select_ln96_4_fu_427_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            dist_fu_64 <= 64'd0;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_reg_499_pp0_iter2_reg == 1'd0))) begin
            dist_fu_64 <= dist_2_reg_561;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                i_fu_68 <= 3'd0;
            end else if (((icmp_ln96_reg_499 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                i_fu_68 <= add_ln293_fu_281_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            idx_fu_80 <= 31'd1;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_fu_186_p2 == 1'd0))) begin
            idx_fu_80 <= select_ln96_2_fu_214_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                indvar_flatten12_fu_84 <= 35'd0;
            end else if (((icmp_ln96_reg_499 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                indvar_flatten12_fu_84 <= add_ln96_fu_276_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            minDist_fu_76 <= minDist_4;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln96_reg_499_pp0_iter9_reg == 1'd0))) begin
            minDist_fu_76 <= select_ln96_3_fu_421_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            add_ln294_reg_515 <= add_ln294_fu_261_p2;
            d_reg_566 <= grp_fu_1462_p_dout0;
            icmp_ln293_reg_503 <= icmp_ln293_fu_200_p2;
            icmp_ln293_reg_503_pp0_iter1_reg <= icmp_ln293_reg_503;
            icmp_ln293_reg_503_pp0_iter2_reg <= icmp_ln293_reg_503_pp0_iter1_reg;
            icmp_ln293_reg_503_pp0_iter3_reg <= icmp_ln293_reg_503_pp0_iter2_reg;
            icmp_ln293_reg_503_pp0_iter4_reg <= icmp_ln293_reg_503_pp0_iter3_reg;
            icmp_ln293_reg_503_pp0_iter5_reg <= icmp_ln293_reg_503_pp0_iter4_reg;
            icmp_ln293_reg_503_pp0_iter6_reg <= icmp_ln293_reg_503_pp0_iter5_reg;
            icmp_ln293_reg_503_pp0_iter7_reg <= icmp_ln293_reg_503_pp0_iter6_reg;
            icmp_ln293_reg_503_pp0_iter8_reg <= icmp_ln293_reg_503_pp0_iter7_reg;
            icmp_ln293_reg_503_pp0_iter9_reg <= icmp_ln293_reg_503_pp0_iter8_reg;
            icmp_ln96_reg_499 <= icmp_ln96_fu_186_p2;
            icmp_ln96_reg_499_pp0_iter1_reg <= icmp_ln96_reg_499;
            icmp_ln96_reg_499_pp0_iter2_reg <= icmp_ln96_reg_499_pp0_iter1_reg;
            icmp_ln96_reg_499_pp0_iter3_reg <= icmp_ln96_reg_499_pp0_iter2_reg;
            icmp_ln96_reg_499_pp0_iter4_reg <= icmp_ln96_reg_499_pp0_iter3_reg;
            icmp_ln96_reg_499_pp0_iter5_reg <= icmp_ln96_reg_499_pp0_iter4_reg;
            icmp_ln96_reg_499_pp0_iter6_reg <= icmp_ln96_reg_499_pp0_iter5_reg;
            icmp_ln96_reg_499_pp0_iter7_reg <= icmp_ln96_reg_499_pp0_iter6_reg;
            icmp_ln96_reg_499_pp0_iter8_reg <= icmp_ln96_reg_499_pp0_iter7_reg;
            icmp_ln96_reg_499_pp0_iter9_reg <= icmp_ln96_reg_499_pp0_iter8_reg;
            idx_2_reg_489 <= idx_fu_80;
            idx_2_reg_489_pp0_iter1_reg <= idx_2_reg_489;
            idx_2_reg_489_pp0_iter2_reg <= idx_2_reg_489_pp0_iter1_reg;
            idx_2_reg_489_pp0_iter3_reg <= idx_2_reg_489_pp0_iter2_reg;
            idx_2_reg_489_pp0_iter4_reg <= idx_2_reg_489_pp0_iter3_reg;
            idx_2_reg_489_pp0_iter5_reg <= idx_2_reg_489_pp0_iter4_reg;
            idx_2_reg_489_pp0_iter6_reg <= idx_2_reg_489_pp0_iter5_reg;
            idx_2_reg_489_pp0_iter7_reg <= idx_2_reg_489_pp0_iter6_reg;
            idx_2_reg_489_pp0_iter8_reg <= idx_2_reg_489_pp0_iter7_reg;
            idx_2_reg_489_pp0_iter9_reg <= idx_2_reg_489_pp0_iter8_reg;
            indvar_flatten12_load_reg_494 <= indvar_flatten12_fu_84;
            mul_i10_i1_reg_556 <= grp_fu_2533_p_dout0;
            select_ln96_1_reg_551 <= select_ln96_1_fu_300_p3;
            select_ln96_reg_510 <= select_ln96_fu_206_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            and_ln98_1_reg_586 <= and_ln98_1_fu_397_p2;
            bestIdx_1_reg_581 <= bestIdx_fu_72;
            bestIdx_3_reg_591 <= bestIdx_3_fu_403_p3;
            rrtVertices_load_reg_535 <= rrtVertices_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            dist_2_reg_561 <= grp_fu_2529_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            goal_load_reg_530 <= goal_q0;
            minDist_1_reg_573 <= minDist_fu_76;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            sub_i9_i1_reg_540 <= grp_fu_2529_p_dout0;
        end
    end

    always @(*) begin
        if (((icmp_ln96_reg_499 == 1'd1) & (1'b0 == ap_block_pp0_stage7_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_condition_exit_pp0_iter0_stage7 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage7 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (icmp_ln96_reg_499_pp0_iter9_reg == 1'd1))) begin
            ap_condition_exit_pp0_iter9_stage3 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter9_stage3 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (~((ap_loop_exit_ready == 1'b0) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter8_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter7_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter6_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter5_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter4_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter1_reg == 1'b0))) begin
            ap_done_pending_pp0 = 1'b1;
        end else begin
            ap_done_pending_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to8 = 1'b1;
        end else begin
            ap_idle_pp0_0to8 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to9 = 1'b1;
        end else begin
            ap_idle_pp0_1to9 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage7_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_reg_499_pp0_iter2_reg == 1'd0))) begin
            ap_sig_allocacmp_dist_1 = dist_2_reg_561;
        end else begin
            ap_sig_allocacmp_dist_1 = dist_fu_64;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (icmp_ln96_reg_499_pp0_iter9_reg == 1'd1))) begin
            bestIdx_6_out_ap_vld = 1'b1;
        end else begin
            bestIdx_6_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            goal_ce0 = 1'b1;
        end else begin
            goal_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln96_reg_499 == 1'd0) & (1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_133_opcode = 2'd1;
        end else if (((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (icmp_ln96_reg_499_pp0_iter2_reg == 1'd0))) begin
            grp_fu_133_opcode = 2'd0;
        end else begin
            grp_fu_133_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_133_p0 = select_ln96_1_reg_551;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_133_p0 = rrtVertices_load_reg_535;
        end else begin
            grp_fu_133_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_133_p1 = mul_i10_i1_reg_556;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_133_p1 = goal_load_reg_530;
        end else begin
            grp_fu_133_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            rrtVertices_ce0 = 1'b1;
        end else begin
            rrtVertices_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_done_pending_pp0 == 1'b0) & (ap_idle_pp0_1to9 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln293_fu_281_p2 = (select_ln96_reg_510 + 3'd1);

    assign add_ln294_fu_261_p2 = (sub_ln294_fu_246_p2 + zext_ln294_fu_257_p1);

    assign add_ln96_1_fu_194_p2 = (idx_fu_80 + 31'd1);

    assign add_ln96_fu_276_p2 = (indvar_flatten12_load_reg_494 + 35'd1);

    assign and_ln98_1_fu_397_p2 = (grp_fu_1454_p_dout0 & and_ln98_fu_391_p2);

    assign and_ln98_fu_391_p2 = (or_ln98_fu_367_p2 & or_ln98_1_fu_385_p2);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage7;

    assign bestIdx_3_fu_403_p3 = ((and_ln98_1_fu_397_p2[0:0] == 1'b1) ? zext_ln96_fu_318_p1 : bestIdx_fu_72);

    assign bestIdx_6_out = bestIdx_3_fu_403_p3[11:0];

    assign bitcast_ln98_1_fu_338_p1 = minDist_1_reg_573;

    assign bitcast_ln98_fu_321_p1 = d_reg_566;

    assign goal_address0 = zext_ln293_fu_252_p1;

    assign grp_fu_1454_p_ce = 1'b1;

    assign grp_fu_1454_p_din0 = d_reg_566;

    assign grp_fu_1454_p_din1 = minDist_fu_76;

    assign grp_fu_1454_p_opcode = 5'd4;

    assign grp_fu_1462_p_ce = 1'b1;

    assign grp_fu_1462_p_din0 = 64'd0;

    assign grp_fu_1462_p_din1 = ap_sig_allocacmp_dist_1;

    assign grp_fu_2529_p_ce = 1'b1;

    assign grp_fu_2529_p_din0 = grp_fu_133_p0;

    assign grp_fu_2529_p_din1 = grp_fu_133_p1;

    assign grp_fu_2529_p_opcode = grp_fu_133_opcode;

    assign grp_fu_2533_p_ce = 1'b1;

    assign grp_fu_2533_p_din0 = sub_i9_i1_reg_540;

    assign grp_fu_2533_p_din1 = sub_i9_i1_reg_540;

    assign icmp_ln293_fu_200_p2 = ((i_fu_68 == 3'd6) ? 1'b1 : 1'b0);

    assign icmp_ln96_fu_186_p2 = ((indvar_flatten12_fu_84 == sub_ln296_1) ? 1'b1 : 1'b0);

    assign icmp_ln98_1_fu_361_p2 = ((trunc_ln98_fu_334_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln98_2_fu_373_p2 = ((tmp_369_dup_fu_341_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln98_3_fu_379_p2 = ((trunc_ln98_1_fu_351_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln98_fu_355_p2 = ((tmp_368_dup_fu_324_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign minDist_6_fu_416_p3 = ((and_ln98_1_reg_586[0:0] == 1'b1) ? d_reg_566 : minDist_1_reg_573);

    assign or_ln98_1_fu_385_p2 = (icmp_ln98_3_fu_379_p2 | icmp_ln98_2_fu_373_p2);

    assign or_ln98_fu_367_p2 = (icmp_ln98_fu_355_p2 | icmp_ln98_1_fu_361_p2);

    assign rrtVertices_address0 = zext_ln294_1_fu_272_p1;

    assign select_ln96_1_fu_300_p3 = ((icmp_ln293_reg_503_pp0_iter1_reg[0:0] == 1'b1) ? 64'd0 : ap_sig_allocacmp_dist_1);

    assign select_ln96_2_fu_214_p3 = ((icmp_ln293_fu_200_p2[0:0] == 1'b1) ? add_ln96_1_fu_194_p2 : idx_fu_80);

    assign select_ln96_3_fu_421_p3 = ((icmp_ln293_reg_503_pp0_iter9_reg[0:0] == 1'b1) ? minDist_6_fu_416_p3 : minDist_1_reg_573);

    assign select_ln96_4_fu_427_p3 = ((icmp_ln293_reg_503_pp0_iter9_reg[0:0] == 1'b1) ? bestIdx_3_reg_591 : bestIdx_1_reg_581);

    assign select_ln96_fu_206_p3 = ((icmp_ln293_fu_200_p2[0:0] == 1'b1) ? 3'd0 : i_fu_68);

    assign sub_ln294_fu_246_p2 = (tmp_33_fu_230_p3 - tmp_34_fu_238_p3);

    assign tmp_33_fu_230_p3 = {{trunc_ln294_1_fu_226_p1}, {3'd0}};

    assign tmp_34_fu_238_p3 = {{trunc_ln294_fu_222_p1}, {1'd0}};

    assign tmp_368_dup_fu_324_p4 = {{bitcast_ln98_fu_321_p1[62:52]}};

    assign tmp_369_dup_fu_341_p4 = {{bitcast_ln98_1_fu_338_p1[62:52]}};

    assign trunc_ln294_1_fu_226_p1 = select_ln96_2_fu_214_p3[9:0];

    assign trunc_ln294_fu_222_p1 = select_ln96_2_fu_214_p3[11:0];

    assign trunc_ln98_1_fu_351_p1 = bitcast_ln98_1_fu_338_p1[51:0];

    assign trunc_ln98_fu_334_p1 = bitcast_ln98_fu_321_p1[51:0];

    assign zext_ln293_fu_252_p1 = select_ln96_fu_206_p3;

    assign zext_ln294_1_fu_272_p1 = add_ln294_reg_515;

    assign zext_ln294_fu_257_p1 = select_ln96_fu_206_p3;

    assign zext_ln96_fu_318_p1 = idx_2_reg_489_pp0_iter9_reg;

endmodule  //main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_110
