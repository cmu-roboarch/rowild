/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    p1_address0,
    p1_ce0,
    p1_q0,
    p1_address1,
    p1_ce1,
    p1_q1,
    p1_offset,
    p2_0_0_address0,
    p2_0_0_ce0,
    p2_0_0_q0,
    p2_0_1_address0,
    p2_0_1_ce0,
    p2_0_1_q0,
    p2_0_2_address0,
    p2_0_2_ce0,
    p2_0_2_q0,
    p2_1_0_address0,
    p2_1_0_ce0,
    p2_1_0_q0,
    p2_1_1_address0,
    p2_1_1_ce0,
    p2_1_1_q0,
    p2_1_2_address0,
    p2_1_2_ce0,
    p2_1_2_q0,
    p2_2_0_address0,
    p2_2_0_ce0,
    p2_2_0_q0,
    p2_2_1_address0,
    p2_2_1_ce0,
    p2_2_1_q0,
    p2_2_2_address0,
    p2_2_2_ce0,
    p2_2_2_q0,
    p2_3_0_address0,
    p2_3_0_ce0,
    p2_3_0_q0,
    p2_3_1_address0,
    p2_3_1_ce0,
    p2_3_1_q0,
    p2_3_2_address0,
    p2_3_2_ce0,
    p2_3_2_q0,
    p2_4_0_address0,
    p2_4_0_ce0,
    p2_4_0_q0,
    p2_4_1_address0,
    p2_4_1_ce0,
    p2_4_1_q0,
    p2_4_2_address0,
    p2_4_2_ce0,
    p2_4_2_q0,
    p2_5_0_address0,
    p2_5_0_ce0,
    p2_5_0_q0,
    p2_5_1_address0,
    p2_5_1_ce0,
    p2_5_1_q0,
    p2_5_2_address0,
    p2_5_2_ce0,
    p2_5_2_q0,
    p2_6_0_address0,
    p2_6_0_ce0,
    p2_6_0_q0,
    p2_6_1_address0,
    p2_6_1_ce0,
    p2_6_1_q0,
    p2_6_2_address0,
    p2_6_2_ce0,
    p2_6_2_q0,
    p2_7_0_address0,
    p2_7_0_ce0,
    p2_7_0_q0,
    p2_7_1_address0,
    p2_7_1_ce0,
    p2_7_1_q0,
    p2_7_2_address0,
    p2_7_2_ce0,
    p2_7_2_q0,
    p2_8_0_address0,
    p2_8_0_ce0,
    p2_8_0_q0,
    p2_8_1_address0,
    p2_8_1_ce0,
    p2_8_1_q0,
    p2_8_2_address0,
    p2_8_2_ce0,
    p2_8_2_q0,
    p2_offset,
    axes1_address0,
    axes1_ce0,
    axes1_q0,
    axes1_address1,
    axes1_ce1,
    axes1_q1,
    ap_return
);

    parameter ap_ST_fsm_state1 = 61'd1;
    parameter ap_ST_fsm_state2 = 61'd2;
    parameter ap_ST_fsm_state3 = 61'd4;
    parameter ap_ST_fsm_state4 = 61'd8;
    parameter ap_ST_fsm_state5 = 61'd16;
    parameter ap_ST_fsm_state6 = 61'd32;
    parameter ap_ST_fsm_state7 = 61'd64;
    parameter ap_ST_fsm_state8 = 61'd128;
    parameter ap_ST_fsm_state9 = 61'd256;
    parameter ap_ST_fsm_state10 = 61'd512;
    parameter ap_ST_fsm_state11 = 61'd1024;
    parameter ap_ST_fsm_state12 = 61'd2048;
    parameter ap_ST_fsm_state13 = 61'd4096;
    parameter ap_ST_fsm_state14 = 61'd8192;
    parameter ap_ST_fsm_state15 = 61'd16384;
    parameter ap_ST_fsm_state16 = 61'd32768;
    parameter ap_ST_fsm_state17 = 61'd65536;
    parameter ap_ST_fsm_state18 = 61'd131072;
    parameter ap_ST_fsm_state19 = 61'd262144;
    parameter ap_ST_fsm_state20 = 61'd524288;
    parameter ap_ST_fsm_state21 = 61'd1048576;
    parameter ap_ST_fsm_state22 = 61'd2097152;
    parameter ap_ST_fsm_state23 = 61'd4194304;
    parameter ap_ST_fsm_state24 = 61'd8388608;
    parameter ap_ST_fsm_state25 = 61'd16777216;
    parameter ap_ST_fsm_state26 = 61'd33554432;
    parameter ap_ST_fsm_state27 = 61'd67108864;
    parameter ap_ST_fsm_state28 = 61'd134217728;
    parameter ap_ST_fsm_state29 = 61'd268435456;
    parameter ap_ST_fsm_state30 = 61'd536870912;
    parameter ap_ST_fsm_state31 = 61'd1073741824;
    parameter ap_ST_fsm_state32 = 61'd2147483648;
    parameter ap_ST_fsm_state33 = 61'd4294967296;
    parameter ap_ST_fsm_state34 = 61'd8589934592;
    parameter ap_ST_fsm_state35 = 61'd17179869184;
    parameter ap_ST_fsm_state36 = 61'd34359738368;
    parameter ap_ST_fsm_state37 = 61'd68719476736;
    parameter ap_ST_fsm_state38 = 61'd137438953472;
    parameter ap_ST_fsm_state39 = 61'd274877906944;
    parameter ap_ST_fsm_state40 = 61'd549755813888;
    parameter ap_ST_fsm_state41 = 61'd1099511627776;
    parameter ap_ST_fsm_state42 = 61'd2199023255552;
    parameter ap_ST_fsm_state43 = 61'd4398046511104;
    parameter ap_ST_fsm_state44 = 61'd8796093022208;
    parameter ap_ST_fsm_state45 = 61'd17592186044416;
    parameter ap_ST_fsm_state46 = 61'd35184372088832;
    parameter ap_ST_fsm_state47 = 61'd70368744177664;
    parameter ap_ST_fsm_state48 = 61'd140737488355328;
    parameter ap_ST_fsm_state49 = 61'd281474976710656;
    parameter ap_ST_fsm_state50 = 61'd562949953421312;
    parameter ap_ST_fsm_state51 = 61'd1125899906842624;
    parameter ap_ST_fsm_state52 = 61'd2251799813685248;
    parameter ap_ST_fsm_state53 = 61'd4503599627370496;
    parameter ap_ST_fsm_state54 = 61'd9007199254740992;
    parameter ap_ST_fsm_state55 = 61'd18014398509481984;
    parameter ap_ST_fsm_state56 = 61'd36028797018963968;
    parameter ap_ST_fsm_state57 = 61'd72057594037927936;
    parameter ap_ST_fsm_state58 = 61'd144115188075855872;
    parameter ap_ST_fsm_state59 = 61'd288230376151711744;
    parameter ap_ST_fsm_state60 = 61'd576460752303423488;
    parameter ap_ST_fsm_state61 = 61'd1152921504606846976;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [6:0] p1_address0;
    output p1_ce0;
    input [63:0] p1_q0;
    output [6:0] p1_address1;
    output p1_ce1;
    input [63:0] p1_q1;
    input [1:0] p1_offset;
    output [2:0] p2_0_0_address0;
    output p2_0_0_ce0;
    input [63:0] p2_0_0_q0;
    output [2:0] p2_0_1_address0;
    output p2_0_1_ce0;
    input [63:0] p2_0_1_q0;
    output [2:0] p2_0_2_address0;
    output p2_0_2_ce0;
    input [63:0] p2_0_2_q0;
    output [2:0] p2_1_0_address0;
    output p2_1_0_ce0;
    input [63:0] p2_1_0_q0;
    output [2:0] p2_1_1_address0;
    output p2_1_1_ce0;
    input [63:0] p2_1_1_q0;
    output [2:0] p2_1_2_address0;
    output p2_1_2_ce0;
    input [63:0] p2_1_2_q0;
    output [2:0] p2_2_0_address0;
    output p2_2_0_ce0;
    input [63:0] p2_2_0_q0;
    output [2:0] p2_2_1_address0;
    output p2_2_1_ce0;
    input [63:0] p2_2_1_q0;
    output [2:0] p2_2_2_address0;
    output p2_2_2_ce0;
    input [63:0] p2_2_2_q0;
    output [2:0] p2_3_0_address0;
    output p2_3_0_ce0;
    input [63:0] p2_3_0_q0;
    output [2:0] p2_3_1_address0;
    output p2_3_1_ce0;
    input [63:0] p2_3_1_q0;
    output [2:0] p2_3_2_address0;
    output p2_3_2_ce0;
    input [63:0] p2_3_2_q0;
    output [2:0] p2_4_0_address0;
    output p2_4_0_ce0;
    input [63:0] p2_4_0_q0;
    output [2:0] p2_4_1_address0;
    output p2_4_1_ce0;
    input [63:0] p2_4_1_q0;
    output [2:0] p2_4_2_address0;
    output p2_4_2_ce0;
    input [63:0] p2_4_2_q0;
    output [2:0] p2_5_0_address0;
    output p2_5_0_ce0;
    input [63:0] p2_5_0_q0;
    output [2:0] p2_5_1_address0;
    output p2_5_1_ce0;
    input [63:0] p2_5_1_q0;
    output [2:0] p2_5_2_address0;
    output p2_5_2_ce0;
    input [63:0] p2_5_2_q0;
    output [2:0] p2_6_0_address0;
    output p2_6_0_ce0;
    input [63:0] p2_6_0_q0;
    output [2:0] p2_6_1_address0;
    output p2_6_1_ce0;
    input [63:0] p2_6_1_q0;
    output [2:0] p2_6_2_address0;
    output p2_6_2_ce0;
    input [63:0] p2_6_2_q0;
    output [2:0] p2_7_0_address0;
    output p2_7_0_ce0;
    input [63:0] p2_7_0_q0;
    output [2:0] p2_7_1_address0;
    output p2_7_1_ce0;
    input [63:0] p2_7_1_q0;
    output [2:0] p2_7_2_address0;
    output p2_7_2_ce0;
    input [63:0] p2_7_2_q0;
    output [2:0] p2_8_0_address0;
    output p2_8_0_ce0;
    input [63:0] p2_8_0_q0;
    output [2:0] p2_8_1_address0;
    output p2_8_1_ce0;
    input [63:0] p2_8_1_q0;
    output [2:0] p2_8_2_address0;
    output p2_8_2_ce0;
    input [63:0] p2_8_2_q0;
    input [2:0] p2_offset;
    output [5:0] axes1_address0;
    output axes1_ce0;
    input [63:0] axes1_q0;
    output [5:0] axes1_address1;
    output axes1_ce1;
    input [63:0] axes1_q1;
    output [0:0] ap_return;

    reg ap_idle;
    reg[0:0] ap_return;

    (* fsm_encoding = "none" *) reg   [60:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire    ap_CS_fsm_state61;
    wire   [0:0] grp_pointsOverlap_double_2_fu_128_ap_return;
    reg   [0:0] icmp_ln166_reg_239;
    reg    ap_condition_exit_pp0_iter0_stage60;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    reg   [0:0] merge_reg_116;
    reg    ap_block_state1_pp0_stage0_iter0;
    reg   [1:0] i_13_reg_234;
    wire   [0:0] icmp_ln166_fu_201_p2;
    wire   [1:0] add_ln166_fu_207_p2;
    reg   [1:0] add_ln166_reg_243;
    wire    grp_pointsOverlap_double_2_fu_128_ap_start;
    wire    grp_pointsOverlap_double_2_fu_128_ap_done;
    wire    grp_pointsOverlap_double_2_fu_128_ap_idle;
    wire    grp_pointsOverlap_double_2_fu_128_ap_ready;
    wire   [6:0] grp_pointsOverlap_double_2_fu_128_p1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p1_ce0;
    wire   [6:0] grp_pointsOverlap_double_2_fu_128_p1_address1;
    wire    grp_pointsOverlap_double_2_fu_128_p1_ce1;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_0_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_0_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_0_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_0_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_0_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_0_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_1_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_1_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_1_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_1_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_1_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_1_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_2_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_2_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_2_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_2_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_2_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_2_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_3_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_3_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_3_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_3_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_3_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_3_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_4_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_4_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_4_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_4_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_4_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_4_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_5_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_5_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_5_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_5_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_5_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_5_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_6_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_6_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_6_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_6_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_6_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_6_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_7_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_7_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_7_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_7_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_7_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_7_2_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_8_0_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_8_0_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_8_1_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_8_1_ce0;
    wire   [2:0] grp_pointsOverlap_double_2_fu_128_p2_8_2_address0;
    wire    grp_pointsOverlap_double_2_fu_128_p2_8_2_ce0;
    wire   [5:0] grp_pointsOverlap_double_2_fu_128_axis_address0;
    wire    grp_pointsOverlap_double_2_fu_128_axis_ce0;
    wire   [5:0] grp_pointsOverlap_double_2_fu_128_axis_address1;
    wire    grp_pointsOverlap_double_2_fu_128_axis_ce1;
    reg   [0:0] ap_phi_mux_merge_phi_fu_120_p4;
    reg    grp_pointsOverlap_double_2_fu_128_ap_start_reg;
    reg   [60:0] ap_NS_fsm;
    wire    ap_NS_fsm_state2;
    wire    ap_CS_fsm_state2;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    wire    ap_CS_fsm_state5;
    wire    ap_CS_fsm_state6;
    wire    ap_CS_fsm_state7;
    wire    ap_CS_fsm_state8;
    wire    ap_CS_fsm_state9;
    wire    ap_CS_fsm_state10;
    wire    ap_CS_fsm_state11;
    wire    ap_CS_fsm_state12;
    wire    ap_CS_fsm_state13;
    wire    ap_CS_fsm_state14;
    wire    ap_CS_fsm_state15;
    wire    ap_CS_fsm_state16;
    wire    ap_CS_fsm_state17;
    reg   [1:0] i_fu_100;
    wire    ap_loop_init;
    reg   [1:0] ap_sig_allocacmp_i_13;
    reg   [0:0] ap_return_preg;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 61'd1;
        #0 grp_pointsOverlap_double_2_fu_128_ap_start_reg = 1'b0;
        #0 i_fu_100 = 2'd0;
        #0 ap_return_preg = 1'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_pointsOverlap_double_2 grp_pointsOverlap_double_2_fu_128 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_pointsOverlap_double_2_fu_128_ap_start),
        .ap_done(grp_pointsOverlap_double_2_fu_128_ap_done),
        .ap_idle(grp_pointsOverlap_double_2_fu_128_ap_idle),
        .ap_ready(grp_pointsOverlap_double_2_fu_128_ap_ready),
        .p1_address0(grp_pointsOverlap_double_2_fu_128_p1_address0),
        .p1_ce0(grp_pointsOverlap_double_2_fu_128_p1_ce0),
        .p1_q0(p1_q0),
        .p1_address1(grp_pointsOverlap_double_2_fu_128_p1_address1),
        .p1_ce1(grp_pointsOverlap_double_2_fu_128_p1_ce1),
        .p1_q1(p1_q1),
        .p1_offset(p1_offset),
        .p2_0_0_address0(grp_pointsOverlap_double_2_fu_128_p2_0_0_address0),
        .p2_0_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_0_0_ce0),
        .p2_0_0_q0(p2_0_0_q0),
        .p2_0_1_address0(grp_pointsOverlap_double_2_fu_128_p2_0_1_address0),
        .p2_0_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_0_1_ce0),
        .p2_0_1_q0(p2_0_1_q0),
        .p2_0_2_address0(grp_pointsOverlap_double_2_fu_128_p2_0_2_address0),
        .p2_0_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_0_2_ce0),
        .p2_0_2_q0(p2_0_2_q0),
        .p2_1_0_address0(grp_pointsOverlap_double_2_fu_128_p2_1_0_address0),
        .p2_1_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_1_0_ce0),
        .p2_1_0_q0(p2_1_0_q0),
        .p2_1_1_address0(grp_pointsOverlap_double_2_fu_128_p2_1_1_address0),
        .p2_1_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_1_1_ce0),
        .p2_1_1_q0(p2_1_1_q0),
        .p2_1_2_address0(grp_pointsOverlap_double_2_fu_128_p2_1_2_address0),
        .p2_1_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_1_2_ce0),
        .p2_1_2_q0(p2_1_2_q0),
        .p2_2_0_address0(grp_pointsOverlap_double_2_fu_128_p2_2_0_address0),
        .p2_2_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_2_0_ce0),
        .p2_2_0_q0(p2_2_0_q0),
        .p2_2_1_address0(grp_pointsOverlap_double_2_fu_128_p2_2_1_address0),
        .p2_2_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_2_1_ce0),
        .p2_2_1_q0(p2_2_1_q0),
        .p2_2_2_address0(grp_pointsOverlap_double_2_fu_128_p2_2_2_address0),
        .p2_2_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_2_2_ce0),
        .p2_2_2_q0(p2_2_2_q0),
        .p2_3_0_address0(grp_pointsOverlap_double_2_fu_128_p2_3_0_address0),
        .p2_3_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_3_0_ce0),
        .p2_3_0_q0(p2_3_0_q0),
        .p2_3_1_address0(grp_pointsOverlap_double_2_fu_128_p2_3_1_address0),
        .p2_3_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_3_1_ce0),
        .p2_3_1_q0(p2_3_1_q0),
        .p2_3_2_address0(grp_pointsOverlap_double_2_fu_128_p2_3_2_address0),
        .p2_3_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_3_2_ce0),
        .p2_3_2_q0(p2_3_2_q0),
        .p2_4_0_address0(grp_pointsOverlap_double_2_fu_128_p2_4_0_address0),
        .p2_4_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_4_0_ce0),
        .p2_4_0_q0(p2_4_0_q0),
        .p2_4_1_address0(grp_pointsOverlap_double_2_fu_128_p2_4_1_address0),
        .p2_4_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_4_1_ce0),
        .p2_4_1_q0(p2_4_1_q0),
        .p2_4_2_address0(grp_pointsOverlap_double_2_fu_128_p2_4_2_address0),
        .p2_4_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_4_2_ce0),
        .p2_4_2_q0(p2_4_2_q0),
        .p2_5_0_address0(grp_pointsOverlap_double_2_fu_128_p2_5_0_address0),
        .p2_5_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_5_0_ce0),
        .p2_5_0_q0(p2_5_0_q0),
        .p2_5_1_address0(grp_pointsOverlap_double_2_fu_128_p2_5_1_address0),
        .p2_5_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_5_1_ce0),
        .p2_5_1_q0(p2_5_1_q0),
        .p2_5_2_address0(grp_pointsOverlap_double_2_fu_128_p2_5_2_address0),
        .p2_5_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_5_2_ce0),
        .p2_5_2_q0(p2_5_2_q0),
        .p2_6_0_address0(grp_pointsOverlap_double_2_fu_128_p2_6_0_address0),
        .p2_6_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_6_0_ce0),
        .p2_6_0_q0(p2_6_0_q0),
        .p2_6_1_address0(grp_pointsOverlap_double_2_fu_128_p2_6_1_address0),
        .p2_6_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_6_1_ce0),
        .p2_6_1_q0(p2_6_1_q0),
        .p2_6_2_address0(grp_pointsOverlap_double_2_fu_128_p2_6_2_address0),
        .p2_6_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_6_2_ce0),
        .p2_6_2_q0(p2_6_2_q0),
        .p2_7_0_address0(grp_pointsOverlap_double_2_fu_128_p2_7_0_address0),
        .p2_7_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_7_0_ce0),
        .p2_7_0_q0(p2_7_0_q0),
        .p2_7_1_address0(grp_pointsOverlap_double_2_fu_128_p2_7_1_address0),
        .p2_7_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_7_1_ce0),
        .p2_7_1_q0(p2_7_1_q0),
        .p2_7_2_address0(grp_pointsOverlap_double_2_fu_128_p2_7_2_address0),
        .p2_7_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_7_2_ce0),
        .p2_7_2_q0(p2_7_2_q0),
        .p2_8_0_address0(grp_pointsOverlap_double_2_fu_128_p2_8_0_address0),
        .p2_8_0_ce0(grp_pointsOverlap_double_2_fu_128_p2_8_0_ce0),
        .p2_8_0_q0(p2_8_0_q0),
        .p2_8_1_address0(grp_pointsOverlap_double_2_fu_128_p2_8_1_address0),
        .p2_8_1_ce0(grp_pointsOverlap_double_2_fu_128_p2_8_1_ce0),
        .p2_8_1_q0(p2_8_1_q0),
        .p2_8_2_address0(grp_pointsOverlap_double_2_fu_128_p2_8_2_address0),
        .p2_8_2_ce0(grp_pointsOverlap_double_2_fu_128_p2_8_2_ce0),
        .p2_8_2_q0(p2_8_2_q0),
        .p2_offset(p2_offset),
        .axis_address0(grp_pointsOverlap_double_2_fu_128_axis_address0),
        .axis_ce0(grp_pointsOverlap_double_2_fu_128_axis_ce0),
        .axis_q0(axes1_q0),
        .axis_address1(grp_pointsOverlap_double_2_fu_128_axis_address1),
        .axis_ce1(grp_pointsOverlap_double_2_fu_128_axis_ce1),
        .axis_q1(axes1_q1),
        .axis_offset1(i_13_reg_234),
        .ap_return(grp_pointsOverlap_double_2_fu_128_ap_return)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage60),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready == 1'b1) & (1'b1 == ap_CS_fsm_state61))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg <= 1'd0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state61) & ((icmp_ln166_reg_239 == 1'd1) | (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd0)))) begin
                ap_return_preg <= ap_phi_mux_merge_phi_fu_120_p4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_pointsOverlap_double_2_fu_128_ap_start_reg <= 1'b0;
        end else begin
            if (((icmp_ln166_fu_201_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1) & (1'b1 == ap_NS_fsm_state2))) begin
                grp_pointsOverlap_double_2_fu_128_ap_start_reg <= 1'b1;
            end else if ((grp_pointsOverlap_double_2_fu_128_ap_ready == 1'b1)) begin
                grp_pointsOverlap_double_2_fu_128_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            i_fu_100 <= 2'd0;
        end else if (((icmp_ln166_reg_239 == 1'd0) & (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd1) & (1'b1 == ap_CS_fsm_state61))) begin
            i_fu_100 <= add_ln166_reg_243;
        end
    end

    always @(posedge ap_clk) begin
        if (((icmp_ln166_reg_239 == 1'd0) & (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state61))) begin
            merge_reg_116 <= 1'd0;
        end else if (((icmp_ln166_fu_201_p2 == 1'd1) & (1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            merge_reg_116 <= 1'd1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
            add_ln166_reg_243 <= add_ln166_fu_207_p2;
            i_13_reg_234 <= ap_sig_allocacmp_i_13;
            icmp_ln166_reg_239 <= icmp_ln166_fu_201_p2;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((1'b1 == ap_block_state1_pp0_stage0_iter0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state61) & ((icmp_ln166_reg_239 == 1'd1) | (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd0)))) begin
            ap_condition_exit_pp0_iter0_stage60 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage60 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready == 1'b1) & (1'b1 == ap_CS_fsm_state61))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln166_reg_239 == 1'd0) & (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd0) & (1'b1 == ap_CS_fsm_state61))) begin
            ap_phi_mux_merge_phi_fu_120_p4 = 1'd0;
        end else begin
            ap_phi_mux_merge_phi_fu_120_p4 = merge_reg_116;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state61)) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state61) & ((icmp_ln166_reg_239 == 1'd1) | (grp_pointsOverlap_double_2_fu_128_ap_return == 1'd0)))) begin
            ap_return = ap_phi_mux_merge_phi_fu_120_p4;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_sig_allocacmp_i_13 = 2'd0;
        end else begin
            ap_sig_allocacmp_i_13 = i_fu_100;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((1'b0 == ap_block_state1_pp0_stage0_iter0) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln166_fu_207_p2 = (ap_sig_allocacmp_i_13 + 2'd1);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];

    assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];

    assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state61 = ap_CS_fsm[32'd60];

    assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign ap_NS_fsm_state2 = ap_NS_fsm[32'd1];

    always @(*) begin
        ap_block_state1_pp0_stage0_iter0 = (ap_start_int == 1'b0);
    end

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage60;

    assign axes1_address0 = grp_pointsOverlap_double_2_fu_128_axis_address0;

    assign axes1_address1 = grp_pointsOverlap_double_2_fu_128_axis_address1;

    assign axes1_ce0 = grp_pointsOverlap_double_2_fu_128_axis_ce0;

    assign axes1_ce1 = grp_pointsOverlap_double_2_fu_128_axis_ce1;

    assign grp_pointsOverlap_double_2_fu_128_ap_start = grp_pointsOverlap_double_2_fu_128_ap_start_reg;

    assign icmp_ln166_fu_201_p2 = ((ap_sig_allocacmp_i_13 == 2'd3) ? 1'b1 : 1'b0);

    assign p1_address0 = grp_pointsOverlap_double_2_fu_128_p1_address0;

    assign p1_address1 = grp_pointsOverlap_double_2_fu_128_p1_address1;

    assign p1_ce0 = grp_pointsOverlap_double_2_fu_128_p1_ce0;

    assign p1_ce1 = grp_pointsOverlap_double_2_fu_128_p1_ce1;

    assign p2_0_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_0_0_address0;

    assign p2_0_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_0_0_ce0;

    assign p2_0_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_0_1_address0;

    assign p2_0_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_0_1_ce0;

    assign p2_0_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_0_2_address0;

    assign p2_0_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_0_2_ce0;

    assign p2_1_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_1_0_address0;

    assign p2_1_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_1_0_ce0;

    assign p2_1_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_1_1_address0;

    assign p2_1_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_1_1_ce0;

    assign p2_1_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_1_2_address0;

    assign p2_1_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_1_2_ce0;

    assign p2_2_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_2_0_address0;

    assign p2_2_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_2_0_ce0;

    assign p2_2_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_2_1_address0;

    assign p2_2_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_2_1_ce0;

    assign p2_2_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_2_2_address0;

    assign p2_2_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_2_2_ce0;

    assign p2_3_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_3_0_address0;

    assign p2_3_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_3_0_ce0;

    assign p2_3_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_3_1_address0;

    assign p2_3_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_3_1_ce0;

    assign p2_3_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_3_2_address0;

    assign p2_3_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_3_2_ce0;

    assign p2_4_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_4_0_address0;

    assign p2_4_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_4_0_ce0;

    assign p2_4_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_4_1_address0;

    assign p2_4_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_4_1_ce0;

    assign p2_4_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_4_2_address0;

    assign p2_4_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_4_2_ce0;

    assign p2_5_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_5_0_address0;

    assign p2_5_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_5_0_ce0;

    assign p2_5_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_5_1_address0;

    assign p2_5_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_5_1_ce0;

    assign p2_5_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_5_2_address0;

    assign p2_5_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_5_2_ce0;

    assign p2_6_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_6_0_address0;

    assign p2_6_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_6_0_ce0;

    assign p2_6_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_6_1_address0;

    assign p2_6_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_6_1_ce0;

    assign p2_6_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_6_2_address0;

    assign p2_6_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_6_2_ce0;

    assign p2_7_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_7_0_address0;

    assign p2_7_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_7_0_ce0;

    assign p2_7_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_7_1_address0;

    assign p2_7_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_7_1_ce0;

    assign p2_7_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_7_2_address0;

    assign p2_7_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_7_2_ce0;

    assign p2_8_0_address0 = grp_pointsOverlap_double_2_fu_128_p2_8_0_address0;

    assign p2_8_0_ce0 = grp_pointsOverlap_double_2_fu_128_p2_8_0_ce0;

    assign p2_8_1_address0 = grp_pointsOverlap_double_2_fu_128_p2_8_1_address0;

    assign p2_8_1_ce0 = grp_pointsOverlap_double_2_fu_128_p2_8_1_ce0;

    assign p2_8_2_address0 = grp_pointsOverlap_double_2_fu_128_p2_8_2_address0;

    assign p2_8_2_ce0 = grp_pointsOverlap_double_2_fu_128_p2_8_2_ce0;

endmodule  //main_cuboidCuboidCollision_double_Pipeline_VITIS_LOOP_166_1
