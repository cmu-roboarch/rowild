/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_48_4 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    state_load_5,
    state_load_4,
    state_load_3,
    state_load_2,
    state_load_1,
    state_load,
    mul,
    mul1,
    mul2,
    add3411_out,
    add3411_out_ap_vld,
    p_out,
    p_out_ap_vld,
    add3010_out,
    add3010_out_ap_vld,
    p_out1,
    p_out1_ap_vld,
    add9_out,
    add9_out_ap_vld,
    p_out2,
    p_out2_ap_vld,
    cost_out,
    cost_out_ap_vld,
    grp_fu_242_p_din0,
    grp_fu_242_p_din1,
    grp_fu_242_p_opcode,
    grp_fu_242_p_dout0,
    grp_fu_242_p_ce,
    grp_fu_247_p_din0,
    grp_fu_247_p_din1,
    grp_fu_247_p_dout0,
    grp_fu_247_p_ce,
    grp_fu_252_p_din0,
    grp_fu_252_p_din1,
    grp_fu_252_p_dout0,
    grp_fu_252_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 5'd1;
    parameter ap_ST_fsm_pp0_stage1 = 5'd2;
    parameter ap_ST_fsm_pp0_stage2 = 5'd4;
    parameter ap_ST_fsm_pp0_stage3 = 5'd8;
    parameter ap_ST_fsm_pp0_stage4 = 5'd16;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [31:0] state_load_5;
    input [31:0] state_load_4;
    input [31:0] state_load_3;
    input [31:0] state_load_2;
    input [31:0] state_load_1;
    input [31:0] state_load;
    input [31:0] mul;
    input [31:0] mul1;
    input [31:0] mul2;
    output [31:0] add3411_out;
    output add3411_out_ap_vld;
    output [31:0] p_out;
    output p_out_ap_vld;
    output [31:0] add3010_out;
    output add3010_out_ap_vld;
    output [31:0] p_out1;
    output p_out1_ap_vld;
    output [31:0] add9_out;
    output add9_out_ap_vld;
    output [31:0] p_out2;
    output p_out2_ap_vld;
    output [31:0] cost_out;
    output cost_out_ap_vld;
    output [31:0] grp_fu_242_p_din0;
    output [31:0] grp_fu_242_p_din1;
    output [0:0] grp_fu_242_p_opcode;
    input [31:0] grp_fu_242_p_dout0;
    output grp_fu_242_p_ce;
    output [31:0] grp_fu_247_p_din0;
    output [31:0] grp_fu_247_p_din1;
    input [31:0] grp_fu_247_p_dout0;
    output grp_fu_247_p_ce;
    output [31:0] grp_fu_252_p_din0;
    output [31:0] grp_fu_252_p_din1;
    input [31:0] grp_fu_252_p_dout0;
    output grp_fu_252_p_ce;

    reg ap_idle;
    reg add3411_out_ap_vld;
    reg p_out_ap_vld;
    reg add3010_out_ap_vld;
    reg p_out1_ap_vld;
    reg add9_out_ap_vld;
    reg p_out2_ap_vld;
    reg cost_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [4:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_subdone;
    reg   [0:0] icmp_ln48_reg_469;
    reg    ap_condition_exit_pp0_iter0_stage4;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    reg   [31:0] reg_232;
    wire    ap_block_pp0_stage0_11001;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire   [31:0] grp_fu_207_p2;
    reg   [31:0] reg_236;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire   [0:0] icmp_ln48_fu_285_p2;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter1_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter2_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter3_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter4_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter5_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter6_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter7_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter8_reg;
    reg   [0:0] icmp_ln48_reg_469_pp0_iter9_reg;
    reg   [31:0] p_load_reg_485;
    reg   [31:0] mul4_reg_491;
    wire    ap_block_pp0_stage4_11001;
    reg   [31:0] mul5_reg_496;
    reg   [31:0] mul6_reg_511;
    wire   [31:0] grp_fu_211_p2;
    reg   [31:0] add5_reg_516;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [31:0] add_reg_526;
    reg   [31:0] add1_reg_532;
    reg   [31:0] add2_reg_538;
    reg   [31:0] sub1_reg_544;
    reg   [31:0] sub3_reg_550;
    reg   [31:0] mul7_reg_556;
    reg   [31:0] mul8_reg_561;
    reg   [31:0] mul9_reg_566;
    reg   [31:0] mul9_reg_566_pp0_iter5_reg;
    reg   [31:0] add6_reg_571;
    reg   [31:0] p_x_assign_reg_576;
    wire   [31:0] grp_fu_227_p2;
    reg   [31:0] tmp_reg_581;
    reg    ap_enable_reg_pp0_iter0_reg;
    reg   [3:0] i_fu_68;
    wire   [3:0] i_2_fu_291_p2;
    wire    ap_loop_init;
    wire    ap_block_pp0_stage1;
    reg   [31:0] cost_fu_72;
    reg   [31:0] ap_sig_allocacmp_cost_load;
    wire    ap_block_pp0_stage4;
    reg   [31:0] empty_fu_76;
    reg   [31:0] ap_sig_allocacmp_p_load19;
    reg   [31:0] add9_fu_80;
    reg   [31:0] ap_sig_allocacmp_add9_load;
    wire    ap_block_pp0_stage0;
    reg   [31:0] empty_9_fu_84;
    reg   [31:0] ap_sig_allocacmp_p_load16;
    reg   [31:0] add3010_fu_88;
    reg   [31:0] ap_sig_allocacmp_add3010_load;
    reg   [31:0] empty_10_fu_92;
    reg   [31:0] ap_sig_allocacmp_p_load;
    reg   [31:0] add3411_fu_96;
    reg   [31:0] ap_sig_allocacmp_add3411_load;
    wire    ap_block_pp0_stage2;
    wire    ap_block_pp0_stage4_01001;
    reg   [31:0] grp_fu_203_p0;
    reg   [31:0] grp_fu_203_p1;
    wire    ap_block_pp0_stage3;
    reg   [31:0] grp_fu_207_p0;
    reg   [31:0] grp_fu_207_p1;
    reg   [31:0] grp_fu_211_p0;
    reg   [31:0] grp_fu_211_p1;
    reg   [31:0] grp_fu_217_p0;
    reg   [31:0] grp_fu_217_p1;
    reg   [31:0] grp_fu_222_p0;
    reg   [31:0] grp_fu_222_p1;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage4_00001;
    reg   [1:0] grp_fu_207_opcode;
    reg   [1:0] grp_fu_211_opcode;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg   [4:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to10;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 5'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 i_fu_68 = 4'd0;
        #0 cost_fu_72 = 32'd0;
        #0 empty_fu_76 = 32'd0;
        #0 add9_fu_80 = 32'd0;
        #0 empty_9_fu_84 = 32'd0;
        #0 add3010_fu_88 = 32'd0;
        #0 empty_10_fu_92 = 32'd0;
        #0 add3411_fu_96 = 32'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_faddfsub_32ns_32ns_32_5_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) faddfsub_32ns_32ns_32_5_full_dsp_1_U5 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_207_p0),
        .din1(grp_fu_207_p1),
        .opcode(grp_fu_207_opcode),
        .ce(1'b1),
        .dout(grp_fu_207_p2)
    );

    main_faddfsub_32ns_32ns_32_5_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) faddfsub_32ns_32ns_32_5_full_dsp_1_U6 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_211_p0),
        .din1(grp_fu_211_p1),
        .opcode(grp_fu_211_opcode),
        .ce(1'b1),
        .dout(grp_fu_211_p2)
    );

    main_fsqrt_32ns_32ns_32_16_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(16),
        .din0_WIDTH(32),
        .din1_WIDTH(32),
        .dout_WIDTH(32)
    ) fsqrt_32ns_32ns_32_16_no_dsp_1_U9 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(32'd0),
        .din1(p_x_assign_reg_576),
        .ce(1'b1),
        .dout(grp_fu_227_p2)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage4),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage4_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage4)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage4_subdone) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                add3010_fu_88 <= state_load_3;
            end else if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
                add3010_fu_88 <= add1_reg_532;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            add3411_fu_96 <= state_load_5;
        end else if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            add3411_fu_96 <= add2_reg_538;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                add9_fu_80 <= state_load_1;
            end else if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
                add9_fu_80 <= add_reg_526;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            cost_fu_72 <= 32'd0;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            cost_fu_72 <= reg_232;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            empty_10_fu_92 <= state_load_4;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            empty_10_fu_92 <= add5_reg_516;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            empty_9_fu_84 <= state_load_2;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            empty_9_fu_84 <= reg_236;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            empty_fu_76 <= state_load;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            empty_fu_76 <= reg_232;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            i_fu_68 <= 4'd0;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln48_fu_285_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            i_fu_68 <= i_2_fu_291_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            add1_reg_532 <= grp_fu_207_p2;
            add_reg_526  <= grp_fu_242_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            add2_reg_538 <= grp_fu_242_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            add5_reg_516 <= grp_fu_211_p2;
            mul6_reg_511 <= grp_fu_247_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            add6_reg_571 <= grp_fu_242_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            icmp_ln48_reg_469 <= icmp_ln48_fu_285_p2;
            icmp_ln48_reg_469_pp0_iter1_reg <= icmp_ln48_reg_469;
            icmp_ln48_reg_469_pp0_iter2_reg <= icmp_ln48_reg_469_pp0_iter1_reg;
            icmp_ln48_reg_469_pp0_iter3_reg <= icmp_ln48_reg_469_pp0_iter2_reg;
            icmp_ln48_reg_469_pp0_iter4_reg <= icmp_ln48_reg_469_pp0_iter3_reg;
            icmp_ln48_reg_469_pp0_iter5_reg <= icmp_ln48_reg_469_pp0_iter4_reg;
            icmp_ln48_reg_469_pp0_iter6_reg <= icmp_ln48_reg_469_pp0_iter5_reg;
            icmp_ln48_reg_469_pp0_iter7_reg <= icmp_ln48_reg_469_pp0_iter6_reg;
            icmp_ln48_reg_469_pp0_iter8_reg <= icmp_ln48_reg_469_pp0_iter7_reg;
            icmp_ln48_reg_469_pp0_iter9_reg <= icmp_ln48_reg_469_pp0_iter8_reg;
            mul9_reg_566_pp0_iter5_reg <= mul9_reg_566;
            p_load_reg_485 <= ap_sig_allocacmp_p_load;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul4_reg_491 <= grp_fu_247_p_dout0;
            mul5_reg_496 <= grp_fu_252_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            mul7_reg_556 <= grp_fu_247_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            mul8_reg_561 <= grp_fu_252_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            mul9_reg_566 <= grp_fu_247_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter6 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            p_x_assign_reg_576 <= grp_fu_207_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            reg_232 <= grp_fu_242_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            reg_236 <= grp_fu_207_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            sub1_reg_544 <= grp_fu_211_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            sub3_reg_550 <= grp_fu_211_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            tmp_reg_581 <= grp_fu_227_p2;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            add3010_out_ap_vld = 1'b1;
        end else begin
            add3010_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            add3411_out_ap_vld = 1'b1;
        end else begin
            add3411_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            add9_out_ap_vld = 1'b1;
        end else begin
            add9_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln48_reg_469 == 1'd1) & (1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_condition_exit_pp0_iter0_stage4 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage4 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to10 = 1'b1;
        end else begin
            ap_idle_pp0_1to10 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_add3010_load = add1_reg_532;
        end else begin
            ap_sig_allocacmp_add3010_load = add3010_fu_88;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_sig_allocacmp_add3411_load = add2_reg_538;
        end else begin
            ap_sig_allocacmp_add3411_load = add3411_fu_96;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_add9_load = add_reg_526;
        end else begin
            ap_sig_allocacmp_add9_load = add9_fu_80;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_sig_allocacmp_cost_load = reg_232;
        end else begin
            ap_sig_allocacmp_cost_load = cost_fu_72;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_sig_allocacmp_p_load = add5_reg_516;
        end else begin
            ap_sig_allocacmp_p_load = empty_10_fu_92;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_sig_allocacmp_p_load16 = reg_236;
        end else begin
            ap_sig_allocacmp_p_load16 = empty_9_fu_84;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_sig_allocacmp_p_load19 = reg_232;
        end else begin
            ap_sig_allocacmp_p_load19 = empty_fu_76;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            cost_out_ap_vld = 1'b1;
        end else begin
            cost_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_203_p0 = ap_sig_allocacmp_cost_load;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_203_p0 = mul7_reg_556;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_203_p0 = ap_sig_allocacmp_add3411_load;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_203_p0 = ap_sig_allocacmp_add9_load;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_203_p0 = ap_sig_allocacmp_p_load19;
        end else begin
            grp_fu_203_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_203_p1 = tmp_reg_581;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_203_p1 = mul8_reg_561;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_203_p1 = mul6_reg_511;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_203_p1 = mul4_reg_491;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_203_p1 = mul;
        end else begin
            grp_fu_203_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_207_opcode = 2'd1;
        end else if ((((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln48_fu_285_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((icmp_ln48_reg_469 == 1'd0) & (1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_207_opcode = 2'd0;
        end else begin
            grp_fu_207_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_207_p0 = add6_reg_571;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_207_p0 = 32'd1092616192;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_207_p0 = ap_sig_allocacmp_add3010_load;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_207_p0 = ap_sig_allocacmp_p_load16;
        end else begin
            grp_fu_207_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter5 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_207_p1 = mul9_reg_566_pp0_iter5_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_207_p1 = add1_reg_532;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_207_p1 = mul5_reg_496;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_207_p1 = mul1;
        end else begin
            grp_fu_207_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_211_opcode = 2'd1;
        end else if (((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln48_fu_285_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_211_opcode = 2'd0;
        end else begin
            grp_fu_211_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_211_p0 = 32'd1092616192;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_211_p0 = ap_sig_allocacmp_p_load;
        end else begin
            grp_fu_211_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_211_p1 = add2_reg_538;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_211_p1 = add_reg_526;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_211_p1 = mul2;
        end else begin
            grp_fu_211_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_217_p0 = sub3_reg_550;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_217_p0 = sub1_reg_544;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_217_p0 = p_load_reg_485;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_217_p0 = ap_sig_allocacmp_p_load19;
        end else begin
            grp_fu_217_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_217_p1 = sub3_reg_550;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_217_p1 = sub1_reg_544;
        end else if ((((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_217_p1 = 32'd1036831949;
        end else begin
            grp_fu_217_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_222_p0 = reg_236;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_222_p0 = ap_sig_allocacmp_p_load16;
        end else begin
            grp_fu_222_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_222_p1 = reg_236;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_222_p1 = 32'd1036831949;
        end else begin
            grp_fu_222_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            p_out1_ap_vld = 1'b1;
        end else begin
            p_out1_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            p_out2_ap_vld = 1'b1;
        end else begin
            p_out2_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (icmp_ln48_reg_469_pp0_iter9_reg == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            p_out_ap_vld = 1'b1;
        end else begin
            p_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to10 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add3010_out = add3010_fu_88;

    assign add3411_out = add3411_fu_96;

    assign add9_out = add9_fu_80;

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage4;

    assign cost_out = cost_fu_72;

    assign grp_fu_242_p_ce = 1'b1;

    assign grp_fu_242_p_din0 = grp_fu_203_p0;

    assign grp_fu_242_p_din1 = grp_fu_203_p1;

    assign grp_fu_242_p_opcode = 2'd0;

    assign grp_fu_247_p_ce = 1'b1;

    assign grp_fu_247_p_din0 = grp_fu_217_p0;

    assign grp_fu_247_p_din1 = grp_fu_217_p1;

    assign grp_fu_252_p_ce = 1'b1;

    assign grp_fu_252_p_din0 = grp_fu_222_p0;

    assign grp_fu_252_p_din1 = grp_fu_222_p1;

    assign i_2_fu_291_p2 = (i_fu_68 + 4'd1);

    assign icmp_ln48_fu_285_p2 = ((i_fu_68 == 4'd10) ? 1'b1 : 1'b0);

    assign p_out = empty_10_fu_92;

    assign p_out1 = empty_9_fu_84;

    assign p_out2 = empty_fu_76;

endmodule  //main_main_Pipeline_VITIS_LOOP_48_4
