/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_56_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    l_TLink_0_0_address0,
    l_TLink_0_0_ce0,
    l_TLink_0_0_we0,
    l_TLink_0_0_d0,
    l_TLink_0_1_address0,
    l_TLink_0_1_ce0,
    l_TLink_0_1_we0,
    l_TLink_0_1_d0,
    l_TLink_0_2_address0,
    l_TLink_0_2_ce0,
    l_TLink_0_2_we0,
    l_TLink_0_2_d0,
    l_TLink_0_3_address0,
    l_TLink_0_3_ce0,
    l_TLink_0_3_we0,
    l_TLink_0_3_d0,
    l_TLink_1_0_address0,
    l_TLink_1_0_ce0,
    l_TLink_1_0_we0,
    l_TLink_1_0_d0,
    l_TLink_1_1_address0,
    l_TLink_1_1_ce0,
    l_TLink_1_1_we0,
    l_TLink_1_1_d0,
    l_TLink_1_2_address0,
    l_TLink_1_2_ce0,
    l_TLink_1_2_we0,
    l_TLink_1_2_d0,
    l_TLink_1_3_address0,
    l_TLink_1_3_ce0,
    l_TLink_1_3_we0,
    l_TLink_1_3_d0,
    l_TLink_2_0_address0,
    l_TLink_2_0_ce0,
    l_TLink_2_0_we0,
    l_TLink_2_0_d0,
    l_TLink_2_1_address0,
    l_TLink_2_1_ce0,
    l_TLink_2_1_we0,
    l_TLink_2_1_d0,
    l_TLink_2_2_address0,
    l_TLink_2_2_ce0,
    l_TLink_2_2_we0,
    l_TLink_2_2_d0,
    l_TLink_2_3_address0,
    l_TLink_2_3_ce0,
    l_TLink_2_3_we0,
    l_TLink_2_3_d0,
    l_TLink_3_0_address0,
    l_TLink_3_0_ce0,
    l_TLink_3_0_we0,
    l_TLink_3_0_d0,
    l_TLink_3_1_address0,
    l_TLink_3_1_ce0,
    l_TLink_3_1_we0,
    l_TLink_3_1_d0,
    l_TLink_3_2_address0,
    l_TLink_3_2_ce0,
    l_TLink_3_2_we0,
    l_TLink_3_2_d0,
    l_TLink_3_3_address0,
    l_TLink_3_3_ce0,
    l_TLink_3_3_we0,
    l_TLink_3_3_d0,
    l_TJoint_0_0_address0,
    l_TJoint_0_0_ce0,
    l_TJoint_0_0_we0,
    l_TJoint_0_0_d0,
    l_TCurr_0_0_address0,
    l_TCurr_0_0_ce0,
    l_TCurr_0_0_we0,
    l_TCurr_0_0_d0,
    l_TJoint_0_1_address0,
    l_TJoint_0_1_ce0,
    l_TJoint_0_1_we0,
    l_TJoint_0_1_d0,
    l_TCurr_0_1_address0,
    l_TCurr_0_1_ce0,
    l_TCurr_0_1_we0,
    l_TCurr_0_1_d0,
    l_TJoint_0_2_address0,
    l_TJoint_0_2_ce0,
    l_TJoint_0_2_we0,
    l_TJoint_0_2_d0,
    l_TCurr_0_2_address0,
    l_TCurr_0_2_ce0,
    l_TCurr_0_2_we0,
    l_TCurr_0_2_d0,
    l_TJoint_0_3_address0,
    l_TJoint_0_3_ce0,
    l_TJoint_0_3_we0,
    l_TJoint_0_3_d0,
    l_TCurr_0_3_address0,
    l_TCurr_0_3_ce0,
    l_TCurr_0_3_we0,
    l_TCurr_0_3_d0,
    l_TJoint_1_0_address0,
    l_TJoint_1_0_ce0,
    l_TJoint_1_0_we0,
    l_TJoint_1_0_d0,
    l_TCurr_1_0_address0,
    l_TCurr_1_0_ce0,
    l_TCurr_1_0_we0,
    l_TCurr_1_0_d0,
    l_TJoint_1_1_address0,
    l_TJoint_1_1_ce0,
    l_TJoint_1_1_we0,
    l_TJoint_1_1_d0,
    l_TCurr_1_1_address0,
    l_TCurr_1_1_ce0,
    l_TCurr_1_1_we0,
    l_TCurr_1_1_d0,
    l_TJoint_1_2_address0,
    l_TJoint_1_2_ce0,
    l_TJoint_1_2_we0,
    l_TJoint_1_2_d0,
    l_TCurr_1_2_address0,
    l_TCurr_1_2_ce0,
    l_TCurr_1_2_we0,
    l_TCurr_1_2_d0,
    l_TJoint_1_3_address0,
    l_TJoint_1_3_ce0,
    l_TJoint_1_3_we0,
    l_TJoint_1_3_d0,
    l_TCurr_1_3_address0,
    l_TCurr_1_3_ce0,
    l_TCurr_1_3_we0,
    l_TCurr_1_3_d0,
    l_TJoint_2_0_address0,
    l_TJoint_2_0_ce0,
    l_TJoint_2_0_we0,
    l_TJoint_2_0_d0,
    l_TCurr_2_0_address0,
    l_TCurr_2_0_ce0,
    l_TCurr_2_0_we0,
    l_TCurr_2_0_d0,
    l_TJoint_2_1_address0,
    l_TJoint_2_1_ce0,
    l_TJoint_2_1_we0,
    l_TJoint_2_1_d0,
    l_TCurr_2_1_address0,
    l_TCurr_2_1_ce0,
    l_TCurr_2_1_we0,
    l_TCurr_2_1_d0,
    l_TJoint_2_2_address0,
    l_TJoint_2_2_ce0,
    l_TJoint_2_2_we0,
    l_TJoint_2_2_d0,
    l_TCurr_2_2_address0,
    l_TCurr_2_2_ce0,
    l_TCurr_2_2_we0,
    l_TCurr_2_2_d0,
    l_TJoint_2_3_address0,
    l_TJoint_2_3_ce0,
    l_TJoint_2_3_we0,
    l_TJoint_2_3_d0,
    l_TCurr_2_3_address0,
    l_TCurr_2_3_ce0,
    l_TCurr_2_3_we0,
    l_TCurr_2_3_d0,
    l_TJoint_3_0_address0,
    l_TJoint_3_0_ce0,
    l_TJoint_3_0_we0,
    l_TJoint_3_0_d0,
    l_TCurr_3_0_address0,
    l_TCurr_3_0_ce0,
    l_TCurr_3_0_we0,
    l_TCurr_3_0_d0,
    l_TJoint_3_1_address0,
    l_TJoint_3_1_ce0,
    l_TJoint_3_1_we0,
    l_TJoint_3_1_d0,
    l_TCurr_3_1_address0,
    l_TCurr_3_1_ce0,
    l_TCurr_3_1_we0,
    l_TCurr_3_1_d0,
    l_TJoint_3_2_address0,
    l_TJoint_3_2_ce0,
    l_TJoint_3_2_we0,
    l_TJoint_3_2_d0,
    l_TCurr_3_2_address0,
    l_TCurr_3_2_ce0,
    l_TCurr_3_2_we0,
    l_TCurr_3_2_d0,
    l_TJoint_3_3_address0,
    l_TJoint_3_3_ce0,
    l_TJoint_3_3_we0,
    l_TJoint_3_3_d0,
    l_TCurr_3_3_address0,
    l_TCurr_3_3_ce0,
    l_TCurr_3_3_we0,
    l_TCurr_3_3_d0
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [2:0] l_TLink_0_0_address0;
    output l_TLink_0_0_ce0;
    output l_TLink_0_0_we0;
    output [63:0] l_TLink_0_0_d0;
    output [2:0] l_TLink_0_1_address0;
    output l_TLink_0_1_ce0;
    output l_TLink_0_1_we0;
    output [63:0] l_TLink_0_1_d0;
    output [2:0] l_TLink_0_2_address0;
    output l_TLink_0_2_ce0;
    output l_TLink_0_2_we0;
    output [63:0] l_TLink_0_2_d0;
    output [2:0] l_TLink_0_3_address0;
    output l_TLink_0_3_ce0;
    output l_TLink_0_3_we0;
    output [63:0] l_TLink_0_3_d0;
    output [2:0] l_TLink_1_0_address0;
    output l_TLink_1_0_ce0;
    output l_TLink_1_0_we0;
    output [63:0] l_TLink_1_0_d0;
    output [2:0] l_TLink_1_1_address0;
    output l_TLink_1_1_ce0;
    output l_TLink_1_1_we0;
    output [63:0] l_TLink_1_1_d0;
    output [2:0] l_TLink_1_2_address0;
    output l_TLink_1_2_ce0;
    output l_TLink_1_2_we0;
    output [63:0] l_TLink_1_2_d0;
    output [2:0] l_TLink_1_3_address0;
    output l_TLink_1_3_ce0;
    output l_TLink_1_3_we0;
    output [63:0] l_TLink_1_3_d0;
    output [2:0] l_TLink_2_0_address0;
    output l_TLink_2_0_ce0;
    output l_TLink_2_0_we0;
    output [63:0] l_TLink_2_0_d0;
    output [2:0] l_TLink_2_1_address0;
    output l_TLink_2_1_ce0;
    output l_TLink_2_1_we0;
    output [63:0] l_TLink_2_1_d0;
    output [2:0] l_TLink_2_2_address0;
    output l_TLink_2_2_ce0;
    output l_TLink_2_2_we0;
    output [63:0] l_TLink_2_2_d0;
    output [2:0] l_TLink_2_3_address0;
    output l_TLink_2_3_ce0;
    output l_TLink_2_3_we0;
    output [63:0] l_TLink_2_3_d0;
    output [2:0] l_TLink_3_0_address0;
    output l_TLink_3_0_ce0;
    output l_TLink_3_0_we0;
    output [63:0] l_TLink_3_0_d0;
    output [2:0] l_TLink_3_1_address0;
    output l_TLink_3_1_ce0;
    output l_TLink_3_1_we0;
    output [63:0] l_TLink_3_1_d0;
    output [2:0] l_TLink_3_2_address0;
    output l_TLink_3_2_ce0;
    output l_TLink_3_2_we0;
    output [63:0] l_TLink_3_2_d0;
    output [2:0] l_TLink_3_3_address0;
    output l_TLink_3_3_ce0;
    output l_TLink_3_3_we0;
    output [63:0] l_TLink_3_3_d0;
    output [2:0] l_TJoint_0_0_address0;
    output l_TJoint_0_0_ce0;
    output l_TJoint_0_0_we0;
    output [63:0] l_TJoint_0_0_d0;
    output [2:0] l_TCurr_0_0_address0;
    output l_TCurr_0_0_ce0;
    output l_TCurr_0_0_we0;
    output [63:0] l_TCurr_0_0_d0;
    output [2:0] l_TJoint_0_1_address0;
    output l_TJoint_0_1_ce0;
    output l_TJoint_0_1_we0;
    output [63:0] l_TJoint_0_1_d0;
    output [2:0] l_TCurr_0_1_address0;
    output l_TCurr_0_1_ce0;
    output l_TCurr_0_1_we0;
    output [63:0] l_TCurr_0_1_d0;
    output [2:0] l_TJoint_0_2_address0;
    output l_TJoint_0_2_ce0;
    output l_TJoint_0_2_we0;
    output [63:0] l_TJoint_0_2_d0;
    output [2:0] l_TCurr_0_2_address0;
    output l_TCurr_0_2_ce0;
    output l_TCurr_0_2_we0;
    output [63:0] l_TCurr_0_2_d0;
    output [2:0] l_TJoint_0_3_address0;
    output l_TJoint_0_3_ce0;
    output l_TJoint_0_3_we0;
    output [63:0] l_TJoint_0_3_d0;
    output [2:0] l_TCurr_0_3_address0;
    output l_TCurr_0_3_ce0;
    output l_TCurr_0_3_we0;
    output [63:0] l_TCurr_0_3_d0;
    output [2:0] l_TJoint_1_0_address0;
    output l_TJoint_1_0_ce0;
    output l_TJoint_1_0_we0;
    output [63:0] l_TJoint_1_0_d0;
    output [2:0] l_TCurr_1_0_address0;
    output l_TCurr_1_0_ce0;
    output l_TCurr_1_0_we0;
    output [63:0] l_TCurr_1_0_d0;
    output [2:0] l_TJoint_1_1_address0;
    output l_TJoint_1_1_ce0;
    output l_TJoint_1_1_we0;
    output [63:0] l_TJoint_1_1_d0;
    output [2:0] l_TCurr_1_1_address0;
    output l_TCurr_1_1_ce0;
    output l_TCurr_1_1_we0;
    output [63:0] l_TCurr_1_1_d0;
    output [2:0] l_TJoint_1_2_address0;
    output l_TJoint_1_2_ce0;
    output l_TJoint_1_2_we0;
    output [63:0] l_TJoint_1_2_d0;
    output [2:0] l_TCurr_1_2_address0;
    output l_TCurr_1_2_ce0;
    output l_TCurr_1_2_we0;
    output [63:0] l_TCurr_1_2_d0;
    output [2:0] l_TJoint_1_3_address0;
    output l_TJoint_1_3_ce0;
    output l_TJoint_1_3_we0;
    output [63:0] l_TJoint_1_3_d0;
    output [2:0] l_TCurr_1_3_address0;
    output l_TCurr_1_3_ce0;
    output l_TCurr_1_3_we0;
    output [63:0] l_TCurr_1_3_d0;
    output [2:0] l_TJoint_2_0_address0;
    output l_TJoint_2_0_ce0;
    output l_TJoint_2_0_we0;
    output [63:0] l_TJoint_2_0_d0;
    output [2:0] l_TCurr_2_0_address0;
    output l_TCurr_2_0_ce0;
    output l_TCurr_2_0_we0;
    output [63:0] l_TCurr_2_0_d0;
    output [2:0] l_TJoint_2_1_address0;
    output l_TJoint_2_1_ce0;
    output l_TJoint_2_1_we0;
    output [63:0] l_TJoint_2_1_d0;
    output [2:0] l_TCurr_2_1_address0;
    output l_TCurr_2_1_ce0;
    output l_TCurr_2_1_we0;
    output [63:0] l_TCurr_2_1_d0;
    output [2:0] l_TJoint_2_2_address0;
    output l_TJoint_2_2_ce0;
    output l_TJoint_2_2_we0;
    output [63:0] l_TJoint_2_2_d0;
    output [2:0] l_TCurr_2_2_address0;
    output l_TCurr_2_2_ce0;
    output l_TCurr_2_2_we0;
    output [63:0] l_TCurr_2_2_d0;
    output [2:0] l_TJoint_2_3_address0;
    output l_TJoint_2_3_ce0;
    output l_TJoint_2_3_we0;
    output [63:0] l_TJoint_2_3_d0;
    output [2:0] l_TCurr_2_3_address0;
    output l_TCurr_2_3_ce0;
    output l_TCurr_2_3_we0;
    output [63:0] l_TCurr_2_3_d0;
    output [2:0] l_TJoint_3_0_address0;
    output l_TJoint_3_0_ce0;
    output l_TJoint_3_0_we0;
    output [63:0] l_TJoint_3_0_d0;
    output [2:0] l_TCurr_3_0_address0;
    output l_TCurr_3_0_ce0;
    output l_TCurr_3_0_we0;
    output [63:0] l_TCurr_3_0_d0;
    output [2:0] l_TJoint_3_1_address0;
    output l_TJoint_3_1_ce0;
    output l_TJoint_3_1_we0;
    output [63:0] l_TJoint_3_1_d0;
    output [2:0] l_TCurr_3_1_address0;
    output l_TCurr_3_1_ce0;
    output l_TCurr_3_1_we0;
    output [63:0] l_TCurr_3_1_d0;
    output [2:0] l_TJoint_3_2_address0;
    output l_TJoint_3_2_ce0;
    output l_TJoint_3_2_we0;
    output [63:0] l_TJoint_3_2_d0;
    output [2:0] l_TCurr_3_2_address0;
    output l_TCurr_3_2_ce0;
    output l_TCurr_3_2_we0;
    output [63:0] l_TCurr_3_2_d0;
    output [2:0] l_TJoint_3_3_address0;
    output l_TJoint_3_3_ce0;
    output l_TJoint_3_3_we0;
    output [63:0] l_TJoint_3_3_d0;
    output [2:0] l_TCurr_3_3_address0;
    output l_TCurr_3_3_ce0;
    output l_TCurr_3_3_we0;
    output [63:0] l_TCurr_3_3_d0;

    reg ap_idle;
    reg l_TJoint_0_0_ce0;
    reg l_TJoint_0_0_we0;
    reg l_TCurr_0_0_ce0;
    reg l_TCurr_0_0_we0;
    reg l_TJoint_0_1_ce0;
    reg l_TJoint_0_1_we0;
    reg l_TCurr_0_1_ce0;
    reg l_TCurr_0_1_we0;
    reg l_TJoint_0_2_ce0;
    reg l_TJoint_0_2_we0;
    reg l_TCurr_0_2_ce0;
    reg l_TCurr_0_2_we0;
    reg l_TJoint_0_3_ce0;
    reg l_TJoint_0_3_we0;
    reg l_TCurr_0_3_ce0;
    reg l_TCurr_0_3_we0;
    reg l_TJoint_1_0_ce0;
    reg l_TJoint_1_0_we0;
    reg l_TCurr_1_0_ce0;
    reg l_TCurr_1_0_we0;
    reg l_TJoint_1_1_ce0;
    reg l_TJoint_1_1_we0;
    reg l_TCurr_1_1_ce0;
    reg l_TCurr_1_1_we0;
    reg l_TJoint_1_2_ce0;
    reg l_TJoint_1_2_we0;
    reg l_TCurr_1_2_ce0;
    reg l_TCurr_1_2_we0;
    reg l_TJoint_1_3_ce0;
    reg l_TJoint_1_3_we0;
    reg l_TCurr_1_3_ce0;
    reg l_TCurr_1_3_we0;
    reg l_TJoint_2_0_ce0;
    reg l_TJoint_2_0_we0;
    reg l_TCurr_2_0_ce0;
    reg l_TCurr_2_0_we0;
    reg l_TJoint_2_1_ce0;
    reg l_TJoint_2_1_we0;
    reg l_TCurr_2_1_ce0;
    reg l_TCurr_2_1_we0;
    reg l_TJoint_2_2_ce0;
    reg l_TJoint_2_2_we0;
    reg l_TCurr_2_2_ce0;
    reg l_TCurr_2_2_we0;
    reg l_TJoint_2_3_ce0;
    reg l_TJoint_2_3_we0;
    reg l_TCurr_2_3_ce0;
    reg l_TCurr_2_3_we0;
    reg l_TJoint_3_0_ce0;
    reg l_TJoint_3_0_we0;
    reg l_TCurr_3_0_ce0;
    reg l_TCurr_3_0_we0;
    reg l_TJoint_3_1_ce0;
    reg l_TJoint_3_1_we0;
    reg l_TCurr_3_1_ce0;
    reg l_TCurr_3_1_we0;
    reg l_TJoint_3_2_ce0;
    reg l_TJoint_3_2_we0;
    reg l_TCurr_3_2_ce0;
    reg l_TCurr_3_2_we0;
    reg l_TJoint_3_3_ce0;
    reg l_TJoint_3_3_we0;
    reg l_TCurr_3_3_ce0;
    reg l_TCurr_3_3_we0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_enable_reg_pp0_iter27;
    reg    ap_enable_reg_pp0_iter28;
    reg    ap_enable_reg_pp0_iter29;
    reg    ap_enable_reg_pp0_iter30;
    reg    ap_enable_reg_pp0_iter31;
    reg    ap_enable_reg_pp0_iter32;
    reg    ap_enable_reg_pp0_iter33;
    reg    ap_enable_reg_pp0_iter34;
    reg    ap_enable_reg_pp0_iter35;
    reg    ap_enable_reg_pp0_iter36;
    reg    ap_enable_reg_pp0_iter37;
    reg    ap_enable_reg_pp0_iter38;
    reg    ap_enable_reg_pp0_iter39;
    reg    ap_enable_reg_pp0_iter40;
    reg    ap_enable_reg_pp0_iter41;
    reg    ap_enable_reg_pp0_iter42;
    reg    ap_enable_reg_pp0_iter43;
    reg    ap_enable_reg_pp0_iter44;
    reg    ap_enable_reg_pp0_iter45;
    reg    ap_enable_reg_pp0_iter46;
    reg    ap_enable_reg_pp0_iter47;
    reg    ap_enable_reg_pp0_iter48;
    reg    ap_enable_reg_pp0_iter49;
    reg    ap_enable_reg_pp0_iter50;
    reg    ap_enable_reg_pp0_iter51;
    reg    ap_enable_reg_pp0_iter52;
    reg    ap_enable_reg_pp0_iter53;
    reg    ap_enable_reg_pp0_iter54;
    reg    ap_enable_reg_pp0_iter55;
    reg    ap_enable_reg_pp0_iter56;
    reg    ap_enable_reg_pp0_iter57;
    reg    ap_enable_reg_pp0_iter58;
    reg    ap_enable_reg_pp0_iter59;
    reg    ap_enable_reg_pp0_iter60;
    reg    ap_enable_reg_pp0_iter61;
    reg    ap_enable_reg_pp0_iter62;
    reg    ap_enable_reg_pp0_iter63;
    reg    ap_enable_reg_pp0_iter64;
    reg    ap_enable_reg_pp0_iter65;
    reg    ap_enable_reg_pp0_iter66;
    reg    ap_enable_reg_pp0_iter67;
    reg    ap_enable_reg_pp0_iter68;
    reg    ap_enable_reg_pp0_iter69;
    reg    ap_enable_reg_pp0_iter70;
    reg    ap_enable_reg_pp0_iter71;
    reg    ap_enable_reg_pp0_iter72;
    reg    ap_enable_reg_pp0_iter73;
    reg    ap_enable_reg_pp0_iter74;
    reg    ap_enable_reg_pp0_iter75;
    reg    ap_enable_reg_pp0_iter76;
    reg    ap_enable_reg_pp0_iter77;
    reg    ap_enable_reg_pp0_iter78;
    reg    ap_enable_reg_pp0_iter79;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    wire   [0:0] icmp_ln56_fu_673_p2;
    reg    ap_condition_exit_pp0_iter0_stage0;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire   [2:0] l_rDesc_3_address0;
    reg    l_rDesc_3_ce0;
    wire   [63:0] l_rDesc_3_q0;
    wire   [2:0] l_rDesc_4_address0;
    reg    l_rDesc_4_ce0;
    wire   [63:0] l_rDesc_4_q0;
    wire   [2:0] l_rDesc_5_address0;
    reg    l_rDesc_5_ce0;
    wire   [63:0] l_rDesc_5_q0;
    reg   [2:0] i_8_reg_736;
    wire    ap_block_pp0_stage0_11001;
    reg   [2:0] i_8_reg_736_pp0_iter1_reg;
    reg   [0:0] icmp_ln56_reg_741;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter1_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter2_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter3_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter4_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter5_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter6_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter7_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter8_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter9_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter10_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter11_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter12_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter13_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter14_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter15_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter16_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter17_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter18_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter19_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter20_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter21_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter22_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter23_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter24_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter25_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter26_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter27_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter28_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter29_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter30_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter31_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter32_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter33_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter34_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter35_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter36_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter37_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter38_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter39_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter40_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter41_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter42_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter43_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter44_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter45_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter46_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter47_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter48_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter49_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter50_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter51_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter52_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter53_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter54_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter55_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter56_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter57_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter58_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter59_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter60_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter61_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter62_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter63_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter64_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter65_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter66_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter67_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter68_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter69_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter70_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter71_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter72_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter73_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter74_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter75_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter76_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter77_reg;
    reg   [0:0] icmp_ln56_reg_741_pp0_iter78_reg;
    reg   [63:0] l_rDesc_3_load_reg_760;
    reg   [63:0] l_rDesc_4_load_reg_765;
    reg   [63:0] l_rDesc_5_load_reg_770;
    wire    grp_rpyxyzToH_double_1_fu_625_ap_start;
    wire    grp_rpyxyzToH_double_1_fu_625_ap_done;
    wire    grp_rpyxyzToH_double_1_fu_625_ap_idle;
    wire    grp_rpyxyzToH_double_1_fu_625_ap_ready;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_0_0_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_0_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_0_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_0_0_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_0_1_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_1_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_1_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_0_1_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_0_2_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_2_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_2_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_0_2_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_0_3_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_3_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_0_3_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_0_3_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_1_0_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_0_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_0_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_1_0_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_1_1_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_1_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_1_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_1_1_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_1_2_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_2_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_2_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_1_2_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_1_3_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_3_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_1_3_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_1_3_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_2_0_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_0_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_0_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_2_0_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_2_1_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_1_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_1_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_2_1_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_2_2_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_2_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_2_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_2_2_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_2_3_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_3_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_2_3_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_2_3_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_3_0_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_0_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_0_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_3_0_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_3_1_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_1_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_1_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_3_1_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_3_2_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_2_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_2_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_3_2_d0;
    wire   [2:0] grp_rpyxyzToH_double_1_fu_625_H_3_3_address0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_3_ce0;
    wire    grp_rpyxyzToH_double_1_fu_625_H_3_3_we0;
    wire   [63:0] grp_rpyxyzToH_double_1_fu_625_H_3_3_d0;
    reg    grp_rpyxyzToH_double_1_fu_625_ap_start_reg;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln56_fu_685_p1;
    reg   [2:0] i_fu_134;
    wire   [2:0] add_ln56_fu_679_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_i_8;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg    ap_loop_exit_ready_pp0_iter10_reg;
    reg    ap_loop_exit_ready_pp0_iter11_reg;
    reg    ap_loop_exit_ready_pp0_iter12_reg;
    reg    ap_loop_exit_ready_pp0_iter13_reg;
    reg    ap_loop_exit_ready_pp0_iter14_reg;
    reg    ap_loop_exit_ready_pp0_iter15_reg;
    reg    ap_loop_exit_ready_pp0_iter16_reg;
    reg    ap_loop_exit_ready_pp0_iter17_reg;
    reg    ap_loop_exit_ready_pp0_iter18_reg;
    reg    ap_loop_exit_ready_pp0_iter19_reg;
    reg    ap_loop_exit_ready_pp0_iter20_reg;
    reg    ap_loop_exit_ready_pp0_iter21_reg;
    reg    ap_loop_exit_ready_pp0_iter22_reg;
    reg    ap_loop_exit_ready_pp0_iter23_reg;
    reg    ap_loop_exit_ready_pp0_iter24_reg;
    reg    ap_loop_exit_ready_pp0_iter25_reg;
    reg    ap_loop_exit_ready_pp0_iter26_reg;
    reg    ap_loop_exit_ready_pp0_iter27_reg;
    reg    ap_loop_exit_ready_pp0_iter28_reg;
    reg    ap_loop_exit_ready_pp0_iter29_reg;
    reg    ap_loop_exit_ready_pp0_iter30_reg;
    reg    ap_loop_exit_ready_pp0_iter31_reg;
    reg    ap_loop_exit_ready_pp0_iter32_reg;
    reg    ap_loop_exit_ready_pp0_iter33_reg;
    reg    ap_loop_exit_ready_pp0_iter34_reg;
    reg    ap_loop_exit_ready_pp0_iter35_reg;
    reg    ap_loop_exit_ready_pp0_iter36_reg;
    reg    ap_loop_exit_ready_pp0_iter37_reg;
    reg    ap_loop_exit_ready_pp0_iter38_reg;
    reg    ap_loop_exit_ready_pp0_iter39_reg;
    reg    ap_loop_exit_ready_pp0_iter40_reg;
    reg    ap_loop_exit_ready_pp0_iter41_reg;
    reg    ap_loop_exit_ready_pp0_iter42_reg;
    reg    ap_loop_exit_ready_pp0_iter43_reg;
    reg    ap_loop_exit_ready_pp0_iter44_reg;
    reg    ap_loop_exit_ready_pp0_iter45_reg;
    reg    ap_loop_exit_ready_pp0_iter46_reg;
    reg    ap_loop_exit_ready_pp0_iter47_reg;
    reg    ap_loop_exit_ready_pp0_iter48_reg;
    reg    ap_loop_exit_ready_pp0_iter49_reg;
    reg    ap_loop_exit_ready_pp0_iter50_reg;
    reg    ap_loop_exit_ready_pp0_iter51_reg;
    reg    ap_loop_exit_ready_pp0_iter52_reg;
    reg    ap_loop_exit_ready_pp0_iter53_reg;
    reg    ap_loop_exit_ready_pp0_iter54_reg;
    reg    ap_loop_exit_ready_pp0_iter55_reg;
    reg    ap_loop_exit_ready_pp0_iter56_reg;
    reg    ap_loop_exit_ready_pp0_iter57_reg;
    reg    ap_loop_exit_ready_pp0_iter58_reg;
    reg    ap_loop_exit_ready_pp0_iter59_reg;
    reg    ap_loop_exit_ready_pp0_iter60_reg;
    reg    ap_loop_exit_ready_pp0_iter61_reg;
    reg    ap_loop_exit_ready_pp0_iter62_reg;
    reg    ap_loop_exit_ready_pp0_iter63_reg;
    reg    ap_loop_exit_ready_pp0_iter64_reg;
    reg    ap_loop_exit_ready_pp0_iter65_reg;
    reg    ap_loop_exit_ready_pp0_iter66_reg;
    reg    ap_loop_exit_ready_pp0_iter67_reg;
    reg    ap_loop_exit_ready_pp0_iter68_reg;
    reg    ap_loop_exit_ready_pp0_iter69_reg;
    reg    ap_loop_exit_ready_pp0_iter70_reg;
    reg    ap_loop_exit_ready_pp0_iter71_reg;
    reg    ap_loop_exit_ready_pp0_iter72_reg;
    reg    ap_loop_exit_ready_pp0_iter73_reg;
    reg    ap_loop_exit_ready_pp0_iter74_reg;
    reg    ap_loop_exit_ready_pp0_iter75_reg;
    reg    ap_loop_exit_ready_pp0_iter76_reg;
    reg    ap_loop_exit_ready_pp0_iter77_reg;
    reg    ap_loop_exit_ready_pp0_iter78_reg;
    reg   [0:0] ap_NS_fsm;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter27 = 1'b0;
        #0 ap_enable_reg_pp0_iter28 = 1'b0;
        #0 ap_enable_reg_pp0_iter29 = 1'b0;
        #0 ap_enable_reg_pp0_iter30 = 1'b0;
        #0 ap_enable_reg_pp0_iter31 = 1'b0;
        #0 ap_enable_reg_pp0_iter32 = 1'b0;
        #0 ap_enable_reg_pp0_iter33 = 1'b0;
        #0 ap_enable_reg_pp0_iter34 = 1'b0;
        #0 ap_enable_reg_pp0_iter35 = 1'b0;
        #0 ap_enable_reg_pp0_iter36 = 1'b0;
        #0 ap_enable_reg_pp0_iter37 = 1'b0;
        #0 ap_enable_reg_pp0_iter38 = 1'b0;
        #0 ap_enable_reg_pp0_iter39 = 1'b0;
        #0 ap_enable_reg_pp0_iter40 = 1'b0;
        #0 ap_enable_reg_pp0_iter41 = 1'b0;
        #0 ap_enable_reg_pp0_iter42 = 1'b0;
        #0 ap_enable_reg_pp0_iter43 = 1'b0;
        #0 ap_enable_reg_pp0_iter44 = 1'b0;
        #0 ap_enable_reg_pp0_iter45 = 1'b0;
        #0 ap_enable_reg_pp0_iter46 = 1'b0;
        #0 ap_enable_reg_pp0_iter47 = 1'b0;
        #0 ap_enable_reg_pp0_iter48 = 1'b0;
        #0 ap_enable_reg_pp0_iter49 = 1'b0;
        #0 ap_enable_reg_pp0_iter50 = 1'b0;
        #0 ap_enable_reg_pp0_iter51 = 1'b0;
        #0 ap_enable_reg_pp0_iter52 = 1'b0;
        #0 ap_enable_reg_pp0_iter53 = 1'b0;
        #0 ap_enable_reg_pp0_iter54 = 1'b0;
        #0 ap_enable_reg_pp0_iter55 = 1'b0;
        #0 ap_enable_reg_pp0_iter56 = 1'b0;
        #0 ap_enable_reg_pp0_iter57 = 1'b0;
        #0 ap_enable_reg_pp0_iter58 = 1'b0;
        #0 ap_enable_reg_pp0_iter59 = 1'b0;
        #0 ap_enable_reg_pp0_iter60 = 1'b0;
        #0 ap_enable_reg_pp0_iter61 = 1'b0;
        #0 ap_enable_reg_pp0_iter62 = 1'b0;
        #0 ap_enable_reg_pp0_iter63 = 1'b0;
        #0 ap_enable_reg_pp0_iter64 = 1'b0;
        #0 ap_enable_reg_pp0_iter65 = 1'b0;
        #0 ap_enable_reg_pp0_iter66 = 1'b0;
        #0 ap_enable_reg_pp0_iter67 = 1'b0;
        #0 ap_enable_reg_pp0_iter68 = 1'b0;
        #0 ap_enable_reg_pp0_iter69 = 1'b0;
        #0 ap_enable_reg_pp0_iter70 = 1'b0;
        #0 ap_enable_reg_pp0_iter71 = 1'b0;
        #0 ap_enable_reg_pp0_iter72 = 1'b0;
        #0 ap_enable_reg_pp0_iter73 = 1'b0;
        #0 ap_enable_reg_pp0_iter74 = 1'b0;
        #0 ap_enable_reg_pp0_iter75 = 1'b0;
        #0 ap_enable_reg_pp0_iter76 = 1'b0;
        #0 ap_enable_reg_pp0_iter77 = 1'b0;
        #0 ap_enable_reg_pp0_iter78 = 1'b0;
        #0 ap_enable_reg_pp0_iter79 = 1'b0;
        #0 grp_rpyxyzToH_double_1_fu_625_ap_start_reg = 1'b0;
        #0 i_fu_134 = 3'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_main_Pipeline_VITIS_LOOP_56_1_l_rDesc_3_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_rDesc_3_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_rDesc_3_address0),
        .ce0(l_rDesc_3_ce0),
        .q0(l_rDesc_3_q0)
    );

    main_main_Pipeline_VITIS_LOOP_56_1_l_rDesc_4_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_rDesc_4_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_rDesc_4_address0),
        .ce0(l_rDesc_4_ce0),
        .q0(l_rDesc_4_q0)
    );

    main_main_Pipeline_VITIS_LOOP_56_1_l_rDesc_5_ROM_AUTO_1R #(
        .DataWidth(64),
        .AddressRange(6),
        .AddressWidth(3)
    ) l_rDesc_5_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(l_rDesc_5_address0),
        .ce0(l_rDesc_5_ce0),
        .q0(l_rDesc_5_q0)
    );

    main_rpyxyzToH_double_1 grp_rpyxyzToH_double_1_fu_625 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_rpyxyzToH_double_1_fu_625_ap_start),
        .ap_done(grp_rpyxyzToH_double_1_fu_625_ap_done),
        .ap_idle(grp_rpyxyzToH_double_1_fu_625_ap_idle),
        .ap_ready(grp_rpyxyzToH_double_1_fu_625_ap_ready),
        .x(l_rDesc_3_load_reg_760),
        .y(l_rDesc_4_load_reg_765),
        .z(l_rDesc_5_load_reg_770),
        .H_0_0_address0(grp_rpyxyzToH_double_1_fu_625_H_0_0_address0),
        .H_0_0_ce0(grp_rpyxyzToH_double_1_fu_625_H_0_0_ce0),
        .H_0_0_we0(grp_rpyxyzToH_double_1_fu_625_H_0_0_we0),
        .H_0_0_d0(grp_rpyxyzToH_double_1_fu_625_H_0_0_d0),
        .H_0_1_address0(grp_rpyxyzToH_double_1_fu_625_H_0_1_address0),
        .H_0_1_ce0(grp_rpyxyzToH_double_1_fu_625_H_0_1_ce0),
        .H_0_1_we0(grp_rpyxyzToH_double_1_fu_625_H_0_1_we0),
        .H_0_1_d0(grp_rpyxyzToH_double_1_fu_625_H_0_1_d0),
        .H_0_2_address0(grp_rpyxyzToH_double_1_fu_625_H_0_2_address0),
        .H_0_2_ce0(grp_rpyxyzToH_double_1_fu_625_H_0_2_ce0),
        .H_0_2_we0(grp_rpyxyzToH_double_1_fu_625_H_0_2_we0),
        .H_0_2_d0(grp_rpyxyzToH_double_1_fu_625_H_0_2_d0),
        .H_0_3_address0(grp_rpyxyzToH_double_1_fu_625_H_0_3_address0),
        .H_0_3_ce0(grp_rpyxyzToH_double_1_fu_625_H_0_3_ce0),
        .H_0_3_we0(grp_rpyxyzToH_double_1_fu_625_H_0_3_we0),
        .H_0_3_d0(grp_rpyxyzToH_double_1_fu_625_H_0_3_d0),
        .H_1_0_address0(grp_rpyxyzToH_double_1_fu_625_H_1_0_address0),
        .H_1_0_ce0(grp_rpyxyzToH_double_1_fu_625_H_1_0_ce0),
        .H_1_0_we0(grp_rpyxyzToH_double_1_fu_625_H_1_0_we0),
        .H_1_0_d0(grp_rpyxyzToH_double_1_fu_625_H_1_0_d0),
        .H_1_1_address0(grp_rpyxyzToH_double_1_fu_625_H_1_1_address0),
        .H_1_1_ce0(grp_rpyxyzToH_double_1_fu_625_H_1_1_ce0),
        .H_1_1_we0(grp_rpyxyzToH_double_1_fu_625_H_1_1_we0),
        .H_1_1_d0(grp_rpyxyzToH_double_1_fu_625_H_1_1_d0),
        .H_1_2_address0(grp_rpyxyzToH_double_1_fu_625_H_1_2_address0),
        .H_1_2_ce0(grp_rpyxyzToH_double_1_fu_625_H_1_2_ce0),
        .H_1_2_we0(grp_rpyxyzToH_double_1_fu_625_H_1_2_we0),
        .H_1_2_d0(grp_rpyxyzToH_double_1_fu_625_H_1_2_d0),
        .H_1_3_address0(grp_rpyxyzToH_double_1_fu_625_H_1_3_address0),
        .H_1_3_ce0(grp_rpyxyzToH_double_1_fu_625_H_1_3_ce0),
        .H_1_3_we0(grp_rpyxyzToH_double_1_fu_625_H_1_3_we0),
        .H_1_3_d0(grp_rpyxyzToH_double_1_fu_625_H_1_3_d0),
        .H_2_0_address0(grp_rpyxyzToH_double_1_fu_625_H_2_0_address0),
        .H_2_0_ce0(grp_rpyxyzToH_double_1_fu_625_H_2_0_ce0),
        .H_2_0_we0(grp_rpyxyzToH_double_1_fu_625_H_2_0_we0),
        .H_2_0_d0(grp_rpyxyzToH_double_1_fu_625_H_2_0_d0),
        .H_2_1_address0(grp_rpyxyzToH_double_1_fu_625_H_2_1_address0),
        .H_2_1_ce0(grp_rpyxyzToH_double_1_fu_625_H_2_1_ce0),
        .H_2_1_we0(grp_rpyxyzToH_double_1_fu_625_H_2_1_we0),
        .H_2_1_d0(grp_rpyxyzToH_double_1_fu_625_H_2_1_d0),
        .H_2_2_address0(grp_rpyxyzToH_double_1_fu_625_H_2_2_address0),
        .H_2_2_ce0(grp_rpyxyzToH_double_1_fu_625_H_2_2_ce0),
        .H_2_2_we0(grp_rpyxyzToH_double_1_fu_625_H_2_2_we0),
        .H_2_2_d0(grp_rpyxyzToH_double_1_fu_625_H_2_2_d0),
        .H_2_3_address0(grp_rpyxyzToH_double_1_fu_625_H_2_3_address0),
        .H_2_3_ce0(grp_rpyxyzToH_double_1_fu_625_H_2_3_ce0),
        .H_2_3_we0(grp_rpyxyzToH_double_1_fu_625_H_2_3_we0),
        .H_2_3_d0(grp_rpyxyzToH_double_1_fu_625_H_2_3_d0),
        .H_3_0_address0(grp_rpyxyzToH_double_1_fu_625_H_3_0_address0),
        .H_3_0_ce0(grp_rpyxyzToH_double_1_fu_625_H_3_0_ce0),
        .H_3_0_we0(grp_rpyxyzToH_double_1_fu_625_H_3_0_we0),
        .H_3_0_d0(grp_rpyxyzToH_double_1_fu_625_H_3_0_d0),
        .H_3_1_address0(grp_rpyxyzToH_double_1_fu_625_H_3_1_address0),
        .H_3_1_ce0(grp_rpyxyzToH_double_1_fu_625_H_3_1_ce0),
        .H_3_1_we0(grp_rpyxyzToH_double_1_fu_625_H_3_1_we0),
        .H_3_1_d0(grp_rpyxyzToH_double_1_fu_625_H_3_1_d0),
        .H_3_2_address0(grp_rpyxyzToH_double_1_fu_625_H_3_2_address0),
        .H_3_2_ce0(grp_rpyxyzToH_double_1_fu_625_H_3_2_ce0),
        .H_3_2_we0(grp_rpyxyzToH_double_1_fu_625_H_3_2_we0),
        .H_3_2_d0(grp_rpyxyzToH_double_1_fu_625_H_3_2_d0),
        .H_3_3_address0(grp_rpyxyzToH_double_1_fu_625_H_3_3_address0),
        .H_3_3_ce0(grp_rpyxyzToH_double_1_fu_625_H_3_3_ce0),
        .H_3_3_we0(grp_rpyxyzToH_double_1_fu_625_H_3_3_we0),
        .H_3_3_d0(grp_rpyxyzToH_double_1_fu_625_H_3_3_d0),
        .H_offset(i_8_reg_736_pp0_iter1_reg)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage0),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready_pp0_iter78_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage0)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter27 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter28 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter29 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter30 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter31 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter32 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter33 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter33 <= ap_enable_reg_pp0_iter32;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter34 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter34 <= ap_enable_reg_pp0_iter33;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter35 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter35 <= ap_enable_reg_pp0_iter34;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter36 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter36 <= ap_enable_reg_pp0_iter35;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter37 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter37 <= ap_enable_reg_pp0_iter36;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter38 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter38 <= ap_enable_reg_pp0_iter37;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter39 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter39 <= ap_enable_reg_pp0_iter38;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter40 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter40 <= ap_enable_reg_pp0_iter39;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter41 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter41 <= ap_enable_reg_pp0_iter40;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter42 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter42 <= ap_enable_reg_pp0_iter41;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter43 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter43 <= ap_enable_reg_pp0_iter42;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter44 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter44 <= ap_enable_reg_pp0_iter43;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter45 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter45 <= ap_enable_reg_pp0_iter44;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter46 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter46 <= ap_enable_reg_pp0_iter45;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter47 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter47 <= ap_enable_reg_pp0_iter46;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter48 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter48 <= ap_enable_reg_pp0_iter47;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter49 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter49 <= ap_enable_reg_pp0_iter48;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter50 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter50 <= ap_enable_reg_pp0_iter49;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter51 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter51 <= ap_enable_reg_pp0_iter50;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter52 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter52 <= ap_enable_reg_pp0_iter51;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter53 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter53 <= ap_enable_reg_pp0_iter52;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter54 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter54 <= ap_enable_reg_pp0_iter53;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter55 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter55 <= ap_enable_reg_pp0_iter54;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter56 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter56 <= ap_enable_reg_pp0_iter55;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter57 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter57 <= ap_enable_reg_pp0_iter56;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter58 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter58 <= ap_enable_reg_pp0_iter57;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter59 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter59 <= ap_enable_reg_pp0_iter58;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter60 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter60 <= ap_enable_reg_pp0_iter59;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter61 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter61 <= ap_enable_reg_pp0_iter60;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter62 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter62 <= ap_enable_reg_pp0_iter61;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter63 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter63 <= ap_enable_reg_pp0_iter62;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter64 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter64 <= ap_enable_reg_pp0_iter63;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter65 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter65 <= ap_enable_reg_pp0_iter64;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter66 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter66 <= ap_enable_reg_pp0_iter65;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter67 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter67 <= ap_enable_reg_pp0_iter66;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter68 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter68 <= ap_enable_reg_pp0_iter67;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter69 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter69 <= ap_enable_reg_pp0_iter68;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter70 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter70 <= ap_enable_reg_pp0_iter69;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter71 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter71 <= ap_enable_reg_pp0_iter70;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter72 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter72 <= ap_enable_reg_pp0_iter71;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter73 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter73 <= ap_enable_reg_pp0_iter72;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter74 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter74 <= ap_enable_reg_pp0_iter73;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter75 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter75 <= ap_enable_reg_pp0_iter74;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter76 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter76 <= ap_enable_reg_pp0_iter75;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter77 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter77 <= ap_enable_reg_pp0_iter76;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter78 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter78 <= ap_enable_reg_pp0_iter77;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter79 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter79 <= ap_enable_reg_pp0_iter78;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_rpyxyzToH_double_1_fu_625_ap_start_reg <= 1'b0;
        end else begin
            if (((icmp_ln56_reg_741 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                grp_rpyxyzToH_double_1_fu_625_ap_start_reg <= 1'b1;
            end else if ((grp_rpyxyzToH_double_1_fu_625_ap_ready == 1'b1)) begin
                grp_rpyxyzToH_double_1_fu_625_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((icmp_ln56_fu_673_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                i_fu_134 <= add_ln56_fu_679_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                i_fu_134 <= 3'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
            ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
            ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
            ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
            ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
            ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
            ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
            ap_loop_exit_ready_pp0_iter17_reg <= ap_loop_exit_ready_pp0_iter16_reg;
            ap_loop_exit_ready_pp0_iter18_reg <= ap_loop_exit_ready_pp0_iter17_reg;
            ap_loop_exit_ready_pp0_iter19_reg <= ap_loop_exit_ready_pp0_iter18_reg;
            ap_loop_exit_ready_pp0_iter20_reg <= ap_loop_exit_ready_pp0_iter19_reg;
            ap_loop_exit_ready_pp0_iter21_reg <= ap_loop_exit_ready_pp0_iter20_reg;
            ap_loop_exit_ready_pp0_iter22_reg <= ap_loop_exit_ready_pp0_iter21_reg;
            ap_loop_exit_ready_pp0_iter23_reg <= ap_loop_exit_ready_pp0_iter22_reg;
            ap_loop_exit_ready_pp0_iter24_reg <= ap_loop_exit_ready_pp0_iter23_reg;
            ap_loop_exit_ready_pp0_iter25_reg <= ap_loop_exit_ready_pp0_iter24_reg;
            ap_loop_exit_ready_pp0_iter26_reg <= ap_loop_exit_ready_pp0_iter25_reg;
            ap_loop_exit_ready_pp0_iter27_reg <= ap_loop_exit_ready_pp0_iter26_reg;
            ap_loop_exit_ready_pp0_iter28_reg <= ap_loop_exit_ready_pp0_iter27_reg;
            ap_loop_exit_ready_pp0_iter29_reg <= ap_loop_exit_ready_pp0_iter28_reg;
            ap_loop_exit_ready_pp0_iter30_reg <= ap_loop_exit_ready_pp0_iter29_reg;
            ap_loop_exit_ready_pp0_iter31_reg <= ap_loop_exit_ready_pp0_iter30_reg;
            ap_loop_exit_ready_pp0_iter32_reg <= ap_loop_exit_ready_pp0_iter31_reg;
            ap_loop_exit_ready_pp0_iter33_reg <= ap_loop_exit_ready_pp0_iter32_reg;
            ap_loop_exit_ready_pp0_iter34_reg <= ap_loop_exit_ready_pp0_iter33_reg;
            ap_loop_exit_ready_pp0_iter35_reg <= ap_loop_exit_ready_pp0_iter34_reg;
            ap_loop_exit_ready_pp0_iter36_reg <= ap_loop_exit_ready_pp0_iter35_reg;
            ap_loop_exit_ready_pp0_iter37_reg <= ap_loop_exit_ready_pp0_iter36_reg;
            ap_loop_exit_ready_pp0_iter38_reg <= ap_loop_exit_ready_pp0_iter37_reg;
            ap_loop_exit_ready_pp0_iter39_reg <= ap_loop_exit_ready_pp0_iter38_reg;
            ap_loop_exit_ready_pp0_iter3_reg  <= ap_loop_exit_ready_pp0_iter2_reg;
            ap_loop_exit_ready_pp0_iter40_reg <= ap_loop_exit_ready_pp0_iter39_reg;
            ap_loop_exit_ready_pp0_iter41_reg <= ap_loop_exit_ready_pp0_iter40_reg;
            ap_loop_exit_ready_pp0_iter42_reg <= ap_loop_exit_ready_pp0_iter41_reg;
            ap_loop_exit_ready_pp0_iter43_reg <= ap_loop_exit_ready_pp0_iter42_reg;
            ap_loop_exit_ready_pp0_iter44_reg <= ap_loop_exit_ready_pp0_iter43_reg;
            ap_loop_exit_ready_pp0_iter45_reg <= ap_loop_exit_ready_pp0_iter44_reg;
            ap_loop_exit_ready_pp0_iter46_reg <= ap_loop_exit_ready_pp0_iter45_reg;
            ap_loop_exit_ready_pp0_iter47_reg <= ap_loop_exit_ready_pp0_iter46_reg;
            ap_loop_exit_ready_pp0_iter48_reg <= ap_loop_exit_ready_pp0_iter47_reg;
            ap_loop_exit_ready_pp0_iter49_reg <= ap_loop_exit_ready_pp0_iter48_reg;
            ap_loop_exit_ready_pp0_iter4_reg  <= ap_loop_exit_ready_pp0_iter3_reg;
            ap_loop_exit_ready_pp0_iter50_reg <= ap_loop_exit_ready_pp0_iter49_reg;
            ap_loop_exit_ready_pp0_iter51_reg <= ap_loop_exit_ready_pp0_iter50_reg;
            ap_loop_exit_ready_pp0_iter52_reg <= ap_loop_exit_ready_pp0_iter51_reg;
            ap_loop_exit_ready_pp0_iter53_reg <= ap_loop_exit_ready_pp0_iter52_reg;
            ap_loop_exit_ready_pp0_iter54_reg <= ap_loop_exit_ready_pp0_iter53_reg;
            ap_loop_exit_ready_pp0_iter55_reg <= ap_loop_exit_ready_pp0_iter54_reg;
            ap_loop_exit_ready_pp0_iter56_reg <= ap_loop_exit_ready_pp0_iter55_reg;
            ap_loop_exit_ready_pp0_iter57_reg <= ap_loop_exit_ready_pp0_iter56_reg;
            ap_loop_exit_ready_pp0_iter58_reg <= ap_loop_exit_ready_pp0_iter57_reg;
            ap_loop_exit_ready_pp0_iter59_reg <= ap_loop_exit_ready_pp0_iter58_reg;
            ap_loop_exit_ready_pp0_iter5_reg  <= ap_loop_exit_ready_pp0_iter4_reg;
            ap_loop_exit_ready_pp0_iter60_reg <= ap_loop_exit_ready_pp0_iter59_reg;
            ap_loop_exit_ready_pp0_iter61_reg <= ap_loop_exit_ready_pp0_iter60_reg;
            ap_loop_exit_ready_pp0_iter62_reg <= ap_loop_exit_ready_pp0_iter61_reg;
            ap_loop_exit_ready_pp0_iter63_reg <= ap_loop_exit_ready_pp0_iter62_reg;
            ap_loop_exit_ready_pp0_iter64_reg <= ap_loop_exit_ready_pp0_iter63_reg;
            ap_loop_exit_ready_pp0_iter65_reg <= ap_loop_exit_ready_pp0_iter64_reg;
            ap_loop_exit_ready_pp0_iter66_reg <= ap_loop_exit_ready_pp0_iter65_reg;
            ap_loop_exit_ready_pp0_iter67_reg <= ap_loop_exit_ready_pp0_iter66_reg;
            ap_loop_exit_ready_pp0_iter68_reg <= ap_loop_exit_ready_pp0_iter67_reg;
            ap_loop_exit_ready_pp0_iter69_reg <= ap_loop_exit_ready_pp0_iter68_reg;
            ap_loop_exit_ready_pp0_iter6_reg  <= ap_loop_exit_ready_pp0_iter5_reg;
            ap_loop_exit_ready_pp0_iter70_reg <= ap_loop_exit_ready_pp0_iter69_reg;
            ap_loop_exit_ready_pp0_iter71_reg <= ap_loop_exit_ready_pp0_iter70_reg;
            ap_loop_exit_ready_pp0_iter72_reg <= ap_loop_exit_ready_pp0_iter71_reg;
            ap_loop_exit_ready_pp0_iter73_reg <= ap_loop_exit_ready_pp0_iter72_reg;
            ap_loop_exit_ready_pp0_iter74_reg <= ap_loop_exit_ready_pp0_iter73_reg;
            ap_loop_exit_ready_pp0_iter75_reg <= ap_loop_exit_ready_pp0_iter74_reg;
            ap_loop_exit_ready_pp0_iter76_reg <= ap_loop_exit_ready_pp0_iter75_reg;
            ap_loop_exit_ready_pp0_iter77_reg <= ap_loop_exit_ready_pp0_iter76_reg;
            ap_loop_exit_ready_pp0_iter78_reg <= ap_loop_exit_ready_pp0_iter77_reg;
            ap_loop_exit_ready_pp0_iter7_reg  <= ap_loop_exit_ready_pp0_iter6_reg;
            ap_loop_exit_ready_pp0_iter8_reg  <= ap_loop_exit_ready_pp0_iter7_reg;
            ap_loop_exit_ready_pp0_iter9_reg  <= ap_loop_exit_ready_pp0_iter8_reg;
            icmp_ln56_reg_741_pp0_iter10_reg  <= icmp_ln56_reg_741_pp0_iter9_reg;
            icmp_ln56_reg_741_pp0_iter11_reg  <= icmp_ln56_reg_741_pp0_iter10_reg;
            icmp_ln56_reg_741_pp0_iter12_reg  <= icmp_ln56_reg_741_pp0_iter11_reg;
            icmp_ln56_reg_741_pp0_iter13_reg  <= icmp_ln56_reg_741_pp0_iter12_reg;
            icmp_ln56_reg_741_pp0_iter14_reg  <= icmp_ln56_reg_741_pp0_iter13_reg;
            icmp_ln56_reg_741_pp0_iter15_reg  <= icmp_ln56_reg_741_pp0_iter14_reg;
            icmp_ln56_reg_741_pp0_iter16_reg  <= icmp_ln56_reg_741_pp0_iter15_reg;
            icmp_ln56_reg_741_pp0_iter17_reg  <= icmp_ln56_reg_741_pp0_iter16_reg;
            icmp_ln56_reg_741_pp0_iter18_reg  <= icmp_ln56_reg_741_pp0_iter17_reg;
            icmp_ln56_reg_741_pp0_iter19_reg  <= icmp_ln56_reg_741_pp0_iter18_reg;
            icmp_ln56_reg_741_pp0_iter20_reg  <= icmp_ln56_reg_741_pp0_iter19_reg;
            icmp_ln56_reg_741_pp0_iter21_reg  <= icmp_ln56_reg_741_pp0_iter20_reg;
            icmp_ln56_reg_741_pp0_iter22_reg  <= icmp_ln56_reg_741_pp0_iter21_reg;
            icmp_ln56_reg_741_pp0_iter23_reg  <= icmp_ln56_reg_741_pp0_iter22_reg;
            icmp_ln56_reg_741_pp0_iter24_reg  <= icmp_ln56_reg_741_pp0_iter23_reg;
            icmp_ln56_reg_741_pp0_iter25_reg  <= icmp_ln56_reg_741_pp0_iter24_reg;
            icmp_ln56_reg_741_pp0_iter26_reg  <= icmp_ln56_reg_741_pp0_iter25_reg;
            icmp_ln56_reg_741_pp0_iter27_reg  <= icmp_ln56_reg_741_pp0_iter26_reg;
            icmp_ln56_reg_741_pp0_iter28_reg  <= icmp_ln56_reg_741_pp0_iter27_reg;
            icmp_ln56_reg_741_pp0_iter29_reg  <= icmp_ln56_reg_741_pp0_iter28_reg;
            icmp_ln56_reg_741_pp0_iter2_reg   <= icmp_ln56_reg_741_pp0_iter1_reg;
            icmp_ln56_reg_741_pp0_iter30_reg  <= icmp_ln56_reg_741_pp0_iter29_reg;
            icmp_ln56_reg_741_pp0_iter31_reg  <= icmp_ln56_reg_741_pp0_iter30_reg;
            icmp_ln56_reg_741_pp0_iter32_reg  <= icmp_ln56_reg_741_pp0_iter31_reg;
            icmp_ln56_reg_741_pp0_iter33_reg  <= icmp_ln56_reg_741_pp0_iter32_reg;
            icmp_ln56_reg_741_pp0_iter34_reg  <= icmp_ln56_reg_741_pp0_iter33_reg;
            icmp_ln56_reg_741_pp0_iter35_reg  <= icmp_ln56_reg_741_pp0_iter34_reg;
            icmp_ln56_reg_741_pp0_iter36_reg  <= icmp_ln56_reg_741_pp0_iter35_reg;
            icmp_ln56_reg_741_pp0_iter37_reg  <= icmp_ln56_reg_741_pp0_iter36_reg;
            icmp_ln56_reg_741_pp0_iter38_reg  <= icmp_ln56_reg_741_pp0_iter37_reg;
            icmp_ln56_reg_741_pp0_iter39_reg  <= icmp_ln56_reg_741_pp0_iter38_reg;
            icmp_ln56_reg_741_pp0_iter3_reg   <= icmp_ln56_reg_741_pp0_iter2_reg;
            icmp_ln56_reg_741_pp0_iter40_reg  <= icmp_ln56_reg_741_pp0_iter39_reg;
            icmp_ln56_reg_741_pp0_iter41_reg  <= icmp_ln56_reg_741_pp0_iter40_reg;
            icmp_ln56_reg_741_pp0_iter42_reg  <= icmp_ln56_reg_741_pp0_iter41_reg;
            icmp_ln56_reg_741_pp0_iter43_reg  <= icmp_ln56_reg_741_pp0_iter42_reg;
            icmp_ln56_reg_741_pp0_iter44_reg  <= icmp_ln56_reg_741_pp0_iter43_reg;
            icmp_ln56_reg_741_pp0_iter45_reg  <= icmp_ln56_reg_741_pp0_iter44_reg;
            icmp_ln56_reg_741_pp0_iter46_reg  <= icmp_ln56_reg_741_pp0_iter45_reg;
            icmp_ln56_reg_741_pp0_iter47_reg  <= icmp_ln56_reg_741_pp0_iter46_reg;
            icmp_ln56_reg_741_pp0_iter48_reg  <= icmp_ln56_reg_741_pp0_iter47_reg;
            icmp_ln56_reg_741_pp0_iter49_reg  <= icmp_ln56_reg_741_pp0_iter48_reg;
            icmp_ln56_reg_741_pp0_iter4_reg   <= icmp_ln56_reg_741_pp0_iter3_reg;
            icmp_ln56_reg_741_pp0_iter50_reg  <= icmp_ln56_reg_741_pp0_iter49_reg;
            icmp_ln56_reg_741_pp0_iter51_reg  <= icmp_ln56_reg_741_pp0_iter50_reg;
            icmp_ln56_reg_741_pp0_iter52_reg  <= icmp_ln56_reg_741_pp0_iter51_reg;
            icmp_ln56_reg_741_pp0_iter53_reg  <= icmp_ln56_reg_741_pp0_iter52_reg;
            icmp_ln56_reg_741_pp0_iter54_reg  <= icmp_ln56_reg_741_pp0_iter53_reg;
            icmp_ln56_reg_741_pp0_iter55_reg  <= icmp_ln56_reg_741_pp0_iter54_reg;
            icmp_ln56_reg_741_pp0_iter56_reg  <= icmp_ln56_reg_741_pp0_iter55_reg;
            icmp_ln56_reg_741_pp0_iter57_reg  <= icmp_ln56_reg_741_pp0_iter56_reg;
            icmp_ln56_reg_741_pp0_iter58_reg  <= icmp_ln56_reg_741_pp0_iter57_reg;
            icmp_ln56_reg_741_pp0_iter59_reg  <= icmp_ln56_reg_741_pp0_iter58_reg;
            icmp_ln56_reg_741_pp0_iter5_reg   <= icmp_ln56_reg_741_pp0_iter4_reg;
            icmp_ln56_reg_741_pp0_iter60_reg  <= icmp_ln56_reg_741_pp0_iter59_reg;
            icmp_ln56_reg_741_pp0_iter61_reg  <= icmp_ln56_reg_741_pp0_iter60_reg;
            icmp_ln56_reg_741_pp0_iter62_reg  <= icmp_ln56_reg_741_pp0_iter61_reg;
            icmp_ln56_reg_741_pp0_iter63_reg  <= icmp_ln56_reg_741_pp0_iter62_reg;
            icmp_ln56_reg_741_pp0_iter64_reg  <= icmp_ln56_reg_741_pp0_iter63_reg;
            icmp_ln56_reg_741_pp0_iter65_reg  <= icmp_ln56_reg_741_pp0_iter64_reg;
            icmp_ln56_reg_741_pp0_iter66_reg  <= icmp_ln56_reg_741_pp0_iter65_reg;
            icmp_ln56_reg_741_pp0_iter67_reg  <= icmp_ln56_reg_741_pp0_iter66_reg;
            icmp_ln56_reg_741_pp0_iter68_reg  <= icmp_ln56_reg_741_pp0_iter67_reg;
            icmp_ln56_reg_741_pp0_iter69_reg  <= icmp_ln56_reg_741_pp0_iter68_reg;
            icmp_ln56_reg_741_pp0_iter6_reg   <= icmp_ln56_reg_741_pp0_iter5_reg;
            icmp_ln56_reg_741_pp0_iter70_reg  <= icmp_ln56_reg_741_pp0_iter69_reg;
            icmp_ln56_reg_741_pp0_iter71_reg  <= icmp_ln56_reg_741_pp0_iter70_reg;
            icmp_ln56_reg_741_pp0_iter72_reg  <= icmp_ln56_reg_741_pp0_iter71_reg;
            icmp_ln56_reg_741_pp0_iter73_reg  <= icmp_ln56_reg_741_pp0_iter72_reg;
            icmp_ln56_reg_741_pp0_iter74_reg  <= icmp_ln56_reg_741_pp0_iter73_reg;
            icmp_ln56_reg_741_pp0_iter75_reg  <= icmp_ln56_reg_741_pp0_iter74_reg;
            icmp_ln56_reg_741_pp0_iter76_reg  <= icmp_ln56_reg_741_pp0_iter75_reg;
            icmp_ln56_reg_741_pp0_iter77_reg  <= icmp_ln56_reg_741_pp0_iter76_reg;
            icmp_ln56_reg_741_pp0_iter78_reg  <= icmp_ln56_reg_741_pp0_iter77_reg;
            icmp_ln56_reg_741_pp0_iter7_reg   <= icmp_ln56_reg_741_pp0_iter6_reg;
            icmp_ln56_reg_741_pp0_iter8_reg   <= icmp_ln56_reg_741_pp0_iter7_reg;
            icmp_ln56_reg_741_pp0_iter9_reg   <= icmp_ln56_reg_741_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
            i_8_reg_736 <= ap_sig_allocacmp_i_8;
            i_8_reg_736_pp0_iter1_reg <= i_8_reg_736;
            icmp_ln56_reg_741 <= icmp_ln56_fu_673_p2;
            icmp_ln56_reg_741_pp0_iter1_reg <= icmp_ln56_reg_741;
            l_rDesc_3_load_reg_760 <= l_rDesc_3_q0;
            l_rDesc_4_load_reg_765 <= l_rDesc_4_q0;
            l_rDesc_5_load_reg_770 <= l_rDesc_5_q0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready_pp0_iter78_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter79 == 1'b0) & (ap_enable_reg_pp0_iter78 == 1'b0) & (ap_enable_reg_pp0_iter77 == 1'b0) 
    & (ap_enable_reg_pp0_iter76 == 1'b0) & (ap_enable_reg_pp0_iter75 == 1'b0) & (ap_enable_reg_pp0_iter74 == 1'b0) & (ap_enable_reg_pp0_iter73 == 1'b0) & (ap_enable_reg_pp0_iter72 == 1'b0) & (ap_enable_reg_pp0_iter71 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter70 == 1'b0) & (ap_enable_reg_pp0_iter69 == 1'b0) & (ap_enable_reg_pp0_iter68 == 1'b0) & (ap_enable_reg_pp0_iter67 == 1'b0) & (ap_enable_reg_pp0_iter66 == 1'b0) & (ap_enable_reg_pp0_iter65 == 1'b0) & (ap_enable_reg_pp0_iter64 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter63 == 1'b0) & (ap_enable_reg_pp0_iter62 == 1'b0) & (ap_enable_reg_pp0_iter61 == 1'b0) & (ap_enable_reg_pp0_iter60 == 1'b0) & (ap_enable_reg_pp0_iter59 == 1'b0) & (ap_enable_reg_pp0_iter58 == 1'b0) & (ap_enable_reg_pp0_iter57 == 1'b0) & (ap_enable_reg_pp0_iter56 == 1'b0) & (ap_enable_reg_pp0_iter55 == 1'b0) & (ap_enable_reg_pp0_iter54 == 1'b0) & (ap_enable_reg_pp0_iter53 == 1'b0) & (ap_enable_reg_pp0_iter52 == 1'b0) & (ap_enable_reg_pp0_iter51 
    == 1'b0) & (ap_enable_reg_pp0_iter50 == 1'b0) & (ap_enable_reg_pp0_iter49 == 1'b0) & (ap_enable_reg_pp0_iter48 == 1'b0) & (ap_enable_reg_pp0_iter47 == 1'b0) & (ap_enable_reg_pp0_iter46 == 1'b0) & (ap_enable_reg_pp0_iter45 == 1'b0) & (ap_enable_reg_pp0_iter44 == 1'b0) & (ap_enable_reg_pp0_iter43 == 1'b0) & (ap_enable_reg_pp0_iter42 == 1'b0) & (ap_enable_reg_pp0_iter41 == 1'b0) & (ap_enable_reg_pp0_iter40 == 1'b0) & (ap_enable_reg_pp0_iter39 == 1'b0) & (ap_enable_reg_pp0_iter38 == 1'b0) & (ap_enable_reg_pp0_iter37 == 1'b0) & (ap_enable_reg_pp0_iter36 == 1'b0) & (ap_enable_reg_pp0_iter35 == 1'b0) & (ap_enable_reg_pp0_iter34 == 1'b0) & (ap_enable_reg_pp0_iter33 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_i_8 = 3'd0;
        end else begin
            ap_sig_allocacmp_i_8 = i_fu_134;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_0_ce0 = 1'b1;
        end else begin
            l_TCurr_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_0_we0 = 1'b1;
        end else begin
            l_TCurr_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_1_ce0 = 1'b1;
        end else begin
            l_TCurr_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_1_we0 = 1'b1;
        end else begin
            l_TCurr_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_2_ce0 = 1'b1;
        end else begin
            l_TCurr_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_2_we0 = 1'b1;
        end else begin
            l_TCurr_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_3_ce0 = 1'b1;
        end else begin
            l_TCurr_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_0_3_we0 = 1'b1;
        end else begin
            l_TCurr_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_0_ce0 = 1'b1;
        end else begin
            l_TCurr_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_0_we0 = 1'b1;
        end else begin
            l_TCurr_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_1_ce0 = 1'b1;
        end else begin
            l_TCurr_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_1_we0 = 1'b1;
        end else begin
            l_TCurr_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_2_ce0 = 1'b1;
        end else begin
            l_TCurr_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_2_we0 = 1'b1;
        end else begin
            l_TCurr_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_3_ce0 = 1'b1;
        end else begin
            l_TCurr_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_1_3_we0 = 1'b1;
        end else begin
            l_TCurr_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_0_ce0 = 1'b1;
        end else begin
            l_TCurr_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_0_we0 = 1'b1;
        end else begin
            l_TCurr_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_1_ce0 = 1'b1;
        end else begin
            l_TCurr_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_1_we0 = 1'b1;
        end else begin
            l_TCurr_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_2_ce0 = 1'b1;
        end else begin
            l_TCurr_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_2_we0 = 1'b1;
        end else begin
            l_TCurr_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_3_ce0 = 1'b1;
        end else begin
            l_TCurr_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_2_3_we0 = 1'b1;
        end else begin
            l_TCurr_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_0_ce0 = 1'b1;
        end else begin
            l_TCurr_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_0_we0 = 1'b1;
        end else begin
            l_TCurr_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_1_ce0 = 1'b1;
        end else begin
            l_TCurr_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_1_we0 = 1'b1;
        end else begin
            l_TCurr_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_2_ce0 = 1'b1;
        end else begin
            l_TCurr_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_2_we0 = 1'b1;
        end else begin
            l_TCurr_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_3_ce0 = 1'b1;
        end else begin
            l_TCurr_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TCurr_3_3_we0 = 1'b1;
        end else begin
            l_TCurr_3_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_0_ce0 = 1'b1;
        end else begin
            l_TJoint_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_0_we0 = 1'b1;
        end else begin
            l_TJoint_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_1_ce0 = 1'b1;
        end else begin
            l_TJoint_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_1_we0 = 1'b1;
        end else begin
            l_TJoint_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_2_ce0 = 1'b1;
        end else begin
            l_TJoint_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_2_we0 = 1'b1;
        end else begin
            l_TJoint_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_3_ce0 = 1'b1;
        end else begin
            l_TJoint_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_0_3_we0 = 1'b1;
        end else begin
            l_TJoint_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_0_ce0 = 1'b1;
        end else begin
            l_TJoint_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_0_we0 = 1'b1;
        end else begin
            l_TJoint_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_1_ce0 = 1'b1;
        end else begin
            l_TJoint_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_1_we0 = 1'b1;
        end else begin
            l_TJoint_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_2_ce0 = 1'b1;
        end else begin
            l_TJoint_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_2_we0 = 1'b1;
        end else begin
            l_TJoint_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_3_ce0 = 1'b1;
        end else begin
            l_TJoint_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_1_3_we0 = 1'b1;
        end else begin
            l_TJoint_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_0_ce0 = 1'b1;
        end else begin
            l_TJoint_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_0_we0 = 1'b1;
        end else begin
            l_TJoint_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_1_ce0 = 1'b1;
        end else begin
            l_TJoint_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_1_we0 = 1'b1;
        end else begin
            l_TJoint_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_2_ce0 = 1'b1;
        end else begin
            l_TJoint_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_2_we0 = 1'b1;
        end else begin
            l_TJoint_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_3_ce0 = 1'b1;
        end else begin
            l_TJoint_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_2_3_we0 = 1'b1;
        end else begin
            l_TJoint_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_0_ce0 = 1'b1;
        end else begin
            l_TJoint_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_0_we0 = 1'b1;
        end else begin
            l_TJoint_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_1_ce0 = 1'b1;
        end else begin
            l_TJoint_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_1_we0 = 1'b1;
        end else begin
            l_TJoint_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_2_ce0 = 1'b1;
        end else begin
            l_TJoint_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_2_we0 = 1'b1;
        end else begin
            l_TJoint_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_3_ce0 = 1'b1;
        end else begin
            l_TJoint_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln56_fu_673_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_TJoint_3_3_we0 = 1'b1;
        end else begin
            l_TJoint_3_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_rDesc_3_ce0 = 1'b1;
        end else begin
            l_rDesc_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_rDesc_4_ce0 = 1'b1;
        end else begin
            l_rDesc_4_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            l_rDesc_5_ce0 = 1'b1;
        end else begin
            l_rDesc_5_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln56_fu_679_p2 = (ap_sig_allocacmp_i_8 + 3'd1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start_int;

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage0;

    assign grp_rpyxyzToH_double_1_fu_625_ap_start = grp_rpyxyzToH_double_1_fu_625_ap_start_reg;

    assign icmp_ln56_fu_673_p2 = ((ap_sig_allocacmp_i_8 == 3'd6) ? 1'b1 : 1'b0);

    assign l_TCurr_0_0_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_0_0_d0 = 64'd4607182418800017408;

    assign l_TCurr_0_1_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_0_1_d0 = 64'd0;

    assign l_TCurr_0_2_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_0_2_d0 = 64'd0;

    assign l_TCurr_0_3_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_0_3_d0 = 64'd0;

    assign l_TCurr_1_0_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_1_0_d0 = 64'd0;

    assign l_TCurr_1_1_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_1_1_d0 = 64'd4607182418800017408;

    assign l_TCurr_1_2_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_1_2_d0 = 64'd0;

    assign l_TCurr_1_3_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_1_3_d0 = 64'd0;

    assign l_TCurr_2_0_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_2_0_d0 = 64'd0;

    assign l_TCurr_2_1_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_2_1_d0 = 64'd0;

    assign l_TCurr_2_2_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_2_2_d0 = 64'd4607182418800017408;

    assign l_TCurr_2_3_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_2_3_d0 = 64'd0;

    assign l_TCurr_3_0_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_3_0_d0 = 64'd0;

    assign l_TCurr_3_1_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_3_1_d0 = 64'd0;

    assign l_TCurr_3_2_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_3_2_d0 = 64'd0;

    assign l_TCurr_3_3_address0 = zext_ln56_fu_685_p1;

    assign l_TCurr_3_3_d0 = 64'd4607182418800017408;

    assign l_TJoint_0_0_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_0_0_d0 = 64'd4607182418800017408;

    assign l_TJoint_0_1_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_0_1_d0 = 64'd0;

    assign l_TJoint_0_2_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_0_2_d0 = 64'd0;

    assign l_TJoint_0_3_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_0_3_d0 = 64'd0;

    assign l_TJoint_1_0_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_1_0_d0 = 64'd0;

    assign l_TJoint_1_1_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_1_1_d0 = 64'd4607182418800017408;

    assign l_TJoint_1_2_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_1_2_d0 = 64'd0;

    assign l_TJoint_1_3_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_1_3_d0 = 64'd0;

    assign l_TJoint_2_0_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_2_0_d0 = 64'd0;

    assign l_TJoint_2_1_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_2_1_d0 = 64'd0;

    assign l_TJoint_2_2_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_2_2_d0 = 64'd4607182418800017408;

    assign l_TJoint_2_3_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_2_3_d0 = 64'd0;

    assign l_TJoint_3_0_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_3_0_d0 = 64'd0;

    assign l_TJoint_3_1_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_3_1_d0 = 64'd0;

    assign l_TJoint_3_2_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_3_2_d0 = 64'd0;

    assign l_TJoint_3_3_address0 = zext_ln56_fu_685_p1;

    assign l_TJoint_3_3_d0 = 64'd4607182418800017408;

    assign l_TLink_0_0_address0 = grp_rpyxyzToH_double_1_fu_625_H_0_0_address0;

    assign l_TLink_0_0_ce0 = grp_rpyxyzToH_double_1_fu_625_H_0_0_ce0;

    assign l_TLink_0_0_d0 = grp_rpyxyzToH_double_1_fu_625_H_0_0_d0;

    assign l_TLink_0_0_we0 = grp_rpyxyzToH_double_1_fu_625_H_0_0_we0;

    assign l_TLink_0_1_address0 = grp_rpyxyzToH_double_1_fu_625_H_0_1_address0;

    assign l_TLink_0_1_ce0 = grp_rpyxyzToH_double_1_fu_625_H_0_1_ce0;

    assign l_TLink_0_1_d0 = grp_rpyxyzToH_double_1_fu_625_H_0_1_d0;

    assign l_TLink_0_1_we0 = grp_rpyxyzToH_double_1_fu_625_H_0_1_we0;

    assign l_TLink_0_2_address0 = grp_rpyxyzToH_double_1_fu_625_H_0_2_address0;

    assign l_TLink_0_2_ce0 = grp_rpyxyzToH_double_1_fu_625_H_0_2_ce0;

    assign l_TLink_0_2_d0 = grp_rpyxyzToH_double_1_fu_625_H_0_2_d0;

    assign l_TLink_0_2_we0 = grp_rpyxyzToH_double_1_fu_625_H_0_2_we0;

    assign l_TLink_0_3_address0 = grp_rpyxyzToH_double_1_fu_625_H_0_3_address0;

    assign l_TLink_0_3_ce0 = grp_rpyxyzToH_double_1_fu_625_H_0_3_ce0;

    assign l_TLink_0_3_d0 = grp_rpyxyzToH_double_1_fu_625_H_0_3_d0;

    assign l_TLink_0_3_we0 = grp_rpyxyzToH_double_1_fu_625_H_0_3_we0;

    assign l_TLink_1_0_address0 = grp_rpyxyzToH_double_1_fu_625_H_1_0_address0;

    assign l_TLink_1_0_ce0 = grp_rpyxyzToH_double_1_fu_625_H_1_0_ce0;

    assign l_TLink_1_0_d0 = grp_rpyxyzToH_double_1_fu_625_H_1_0_d0;

    assign l_TLink_1_0_we0 = grp_rpyxyzToH_double_1_fu_625_H_1_0_we0;

    assign l_TLink_1_1_address0 = grp_rpyxyzToH_double_1_fu_625_H_1_1_address0;

    assign l_TLink_1_1_ce0 = grp_rpyxyzToH_double_1_fu_625_H_1_1_ce0;

    assign l_TLink_1_1_d0 = grp_rpyxyzToH_double_1_fu_625_H_1_1_d0;

    assign l_TLink_1_1_we0 = grp_rpyxyzToH_double_1_fu_625_H_1_1_we0;

    assign l_TLink_1_2_address0 = grp_rpyxyzToH_double_1_fu_625_H_1_2_address0;

    assign l_TLink_1_2_ce0 = grp_rpyxyzToH_double_1_fu_625_H_1_2_ce0;

    assign l_TLink_1_2_d0 = grp_rpyxyzToH_double_1_fu_625_H_1_2_d0;

    assign l_TLink_1_2_we0 = grp_rpyxyzToH_double_1_fu_625_H_1_2_we0;

    assign l_TLink_1_3_address0 = grp_rpyxyzToH_double_1_fu_625_H_1_3_address0;

    assign l_TLink_1_3_ce0 = grp_rpyxyzToH_double_1_fu_625_H_1_3_ce0;

    assign l_TLink_1_3_d0 = grp_rpyxyzToH_double_1_fu_625_H_1_3_d0;

    assign l_TLink_1_3_we0 = grp_rpyxyzToH_double_1_fu_625_H_1_3_we0;

    assign l_TLink_2_0_address0 = grp_rpyxyzToH_double_1_fu_625_H_2_0_address0;

    assign l_TLink_2_0_ce0 = grp_rpyxyzToH_double_1_fu_625_H_2_0_ce0;

    assign l_TLink_2_0_d0 = grp_rpyxyzToH_double_1_fu_625_H_2_0_d0;

    assign l_TLink_2_0_we0 = grp_rpyxyzToH_double_1_fu_625_H_2_0_we0;

    assign l_TLink_2_1_address0 = grp_rpyxyzToH_double_1_fu_625_H_2_1_address0;

    assign l_TLink_2_1_ce0 = grp_rpyxyzToH_double_1_fu_625_H_2_1_ce0;

    assign l_TLink_2_1_d0 = grp_rpyxyzToH_double_1_fu_625_H_2_1_d0;

    assign l_TLink_2_1_we0 = grp_rpyxyzToH_double_1_fu_625_H_2_1_we0;

    assign l_TLink_2_2_address0 = grp_rpyxyzToH_double_1_fu_625_H_2_2_address0;

    assign l_TLink_2_2_ce0 = grp_rpyxyzToH_double_1_fu_625_H_2_2_ce0;

    assign l_TLink_2_2_d0 = grp_rpyxyzToH_double_1_fu_625_H_2_2_d0;

    assign l_TLink_2_2_we0 = grp_rpyxyzToH_double_1_fu_625_H_2_2_we0;

    assign l_TLink_2_3_address0 = grp_rpyxyzToH_double_1_fu_625_H_2_3_address0;

    assign l_TLink_2_3_ce0 = grp_rpyxyzToH_double_1_fu_625_H_2_3_ce0;

    assign l_TLink_2_3_d0 = grp_rpyxyzToH_double_1_fu_625_H_2_3_d0;

    assign l_TLink_2_3_we0 = grp_rpyxyzToH_double_1_fu_625_H_2_3_we0;

    assign l_TLink_3_0_address0 = grp_rpyxyzToH_double_1_fu_625_H_3_0_address0;

    assign l_TLink_3_0_ce0 = grp_rpyxyzToH_double_1_fu_625_H_3_0_ce0;

    assign l_TLink_3_0_d0 = grp_rpyxyzToH_double_1_fu_625_H_3_0_d0;

    assign l_TLink_3_0_we0 = grp_rpyxyzToH_double_1_fu_625_H_3_0_we0;

    assign l_TLink_3_1_address0 = grp_rpyxyzToH_double_1_fu_625_H_3_1_address0;

    assign l_TLink_3_1_ce0 = grp_rpyxyzToH_double_1_fu_625_H_3_1_ce0;

    assign l_TLink_3_1_d0 = grp_rpyxyzToH_double_1_fu_625_H_3_1_d0;

    assign l_TLink_3_1_we0 = grp_rpyxyzToH_double_1_fu_625_H_3_1_we0;

    assign l_TLink_3_2_address0 = grp_rpyxyzToH_double_1_fu_625_H_3_2_address0;

    assign l_TLink_3_2_ce0 = grp_rpyxyzToH_double_1_fu_625_H_3_2_ce0;

    assign l_TLink_3_2_d0 = grp_rpyxyzToH_double_1_fu_625_H_3_2_d0;

    assign l_TLink_3_2_we0 = grp_rpyxyzToH_double_1_fu_625_H_3_2_we0;

    assign l_TLink_3_3_address0 = grp_rpyxyzToH_double_1_fu_625_H_3_3_address0;

    assign l_TLink_3_3_ce0 = grp_rpyxyzToH_double_1_fu_625_H_3_3_ce0;

    assign l_TLink_3_3_d0 = grp_rpyxyzToH_double_1_fu_625_H_3_3_d0;

    assign l_TLink_3_3_we0 = grp_rpyxyzToH_double_1_fu_625_H_3_3_we0;

    assign l_rDesc_3_address0 = zext_ln56_fu_685_p1;

    assign l_rDesc_4_address0 = zext_ln56_fu_685_p1;

    assign l_rDesc_5_address0 = zext_ln56_fu_685_p1;

    assign zext_ln56_fu_685_p1 = ap_sig_allocacmp_i_8;

endmodule  //main_main_Pipeline_VITIS_LOOP_56_1
