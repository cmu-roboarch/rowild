/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_rpyxyzToH_double_s (
    ap_clk,
    ap_rst,
    x,
    y,
    z,
    p_read,
    p_read1,
    p_read2,
    p_read3,
    p_read4,
    p_read5,
    p_read6,
    p_read7,
    p_read8,
    p_read9,
    p_read10,
    p_read11,
    p_read12,
    p_read13,
    p_read14,
    p_read15,
    p_read16,
    p_read17,
    p_read18,
    p_read19,
    p_read20,
    p_read21,
    p_read22,
    p_read23,
    p_read24,
    p_read25,
    p_read26,
    p_read27,
    p_read28,
    p_read29,
    p_read30,
    p_read31,
    p_read32,
    p_read33,
    p_read34,
    p_read35,
    p_read36,
    p_read37,
    p_read38,
    p_read39,
    p_read40,
    p_read41,
    p_read42,
    p_read43,
    p_read44,
    p_read45,
    p_read46,
    p_read47,
    p_read48,
    p_read49,
    p_read50,
    p_read51,
    p_read52,
    p_read53,
    p_read54,
    p_read55,
    p_read56,
    p_read57,
    p_read58,
    p_read59,
    p_read60,
    p_read61,
    p_read62,
    p_read63,
    H_offset,
    ap_return_0,
    ap_return_1,
    ap_return_2,
    ap_return_3,
    ap_return_4,
    ap_return_5,
    ap_return_6,
    ap_return_7,
    ap_return_8,
    ap_return_9,
    ap_return_10,
    ap_return_11,
    ap_return_12,
    ap_return_13,
    ap_return_14,
    ap_return_15,
    ap_return_16,
    ap_return_17,
    ap_return_18,
    ap_return_19,
    ap_return_20,
    ap_return_21,
    ap_return_22,
    ap_return_23,
    ap_return_24,
    ap_return_25,
    ap_return_26,
    ap_return_27,
    ap_return_28,
    ap_return_29,
    ap_return_30,
    ap_return_31,
    ap_return_32,
    ap_return_33,
    ap_return_34,
    ap_return_35,
    ap_return_36,
    ap_return_37,
    ap_return_38,
    ap_return_39,
    ap_return_40,
    ap_return_41,
    ap_return_42,
    ap_return_43,
    ap_return_44,
    ap_return_45,
    ap_return_46,
    ap_return_47,
    ap_return_48,
    ap_return_49,
    ap_return_50,
    ap_return_51,
    ap_return_52,
    ap_return_53,
    ap_return_54,
    ap_return_55,
    ap_return_56,
    ap_return_57,
    ap_return_58,
    ap_return_59,
    ap_return_60,
    ap_return_61,
    ap_return_62,
    ap_return_63
);


    input ap_clk;
    input ap_rst;
    input [63:0] x;
    input [63:0] y;
    input [63:0] z;
    input [63:0] p_read;
    input [63:0] p_read1;
    input [63:0] p_read2;
    input [63:0] p_read3;
    input [63:0] p_read4;
    input [63:0] p_read5;
    input [63:0] p_read6;
    input [63:0] p_read7;
    input [63:0] p_read8;
    input [63:0] p_read9;
    input [63:0] p_read10;
    input [63:0] p_read11;
    input [63:0] p_read12;
    input [63:0] p_read13;
    input [63:0] p_read14;
    input [63:0] p_read15;
    input [63:0] p_read16;
    input [63:0] p_read17;
    input [63:0] p_read18;
    input [63:0] p_read19;
    input [63:0] p_read20;
    input [63:0] p_read21;
    input [63:0] p_read22;
    input [63:0] p_read23;
    input [63:0] p_read24;
    input [63:0] p_read25;
    input [63:0] p_read26;
    input [63:0] p_read27;
    input [63:0] p_read28;
    input [63:0] p_read29;
    input [63:0] p_read30;
    input [63:0] p_read31;
    input [63:0] p_read32;
    input [63:0] p_read33;
    input [63:0] p_read34;
    input [63:0] p_read35;
    input [63:0] p_read36;
    input [63:0] p_read37;
    input [63:0] p_read38;
    input [63:0] p_read39;
    input [63:0] p_read40;
    input [63:0] p_read41;
    input [63:0] p_read42;
    input [63:0] p_read43;
    input [63:0] p_read44;
    input [63:0] p_read45;
    input [63:0] p_read46;
    input [63:0] p_read47;
    input [63:0] p_read48;
    input [63:0] p_read49;
    input [63:0] p_read50;
    input [63:0] p_read51;
    input [63:0] p_read52;
    input [63:0] p_read53;
    input [63:0] p_read54;
    input [63:0] p_read55;
    input [63:0] p_read56;
    input [63:0] p_read57;
    input [63:0] p_read58;
    input [63:0] p_read59;
    input [63:0] p_read60;
    input [63:0] p_read61;
    input [63:0] p_read62;
    input [63:0] p_read63;
    input [1:0] H_offset;
    output [63:0] ap_return_0;
    output [63:0] ap_return_1;
    output [63:0] ap_return_2;
    output [63:0] ap_return_3;
    output [63:0] ap_return_4;
    output [63:0] ap_return_5;
    output [63:0] ap_return_6;
    output [63:0] ap_return_7;
    output [63:0] ap_return_8;
    output [63:0] ap_return_9;
    output [63:0] ap_return_10;
    output [63:0] ap_return_11;
    output [63:0] ap_return_12;
    output [63:0] ap_return_13;
    output [63:0] ap_return_14;
    output [63:0] ap_return_15;
    output [63:0] ap_return_16;
    output [63:0] ap_return_17;
    output [63:0] ap_return_18;
    output [63:0] ap_return_19;
    output [63:0] ap_return_20;
    output [63:0] ap_return_21;
    output [63:0] ap_return_22;
    output [63:0] ap_return_23;
    output [63:0] ap_return_24;
    output [63:0] ap_return_25;
    output [63:0] ap_return_26;
    output [63:0] ap_return_27;
    output [63:0] ap_return_28;
    output [63:0] ap_return_29;
    output [63:0] ap_return_30;
    output [63:0] ap_return_31;
    output [63:0] ap_return_32;
    output [63:0] ap_return_33;
    output [63:0] ap_return_34;
    output [63:0] ap_return_35;
    output [63:0] ap_return_36;
    output [63:0] ap_return_37;
    output [63:0] ap_return_38;
    output [63:0] ap_return_39;
    output [63:0] ap_return_40;
    output [63:0] ap_return_41;
    output [63:0] ap_return_42;
    output [63:0] ap_return_43;
    output [63:0] ap_return_44;
    output [63:0] ap_return_45;
    output [63:0] ap_return_46;
    output [63:0] ap_return_47;
    output [63:0] ap_return_48;
    output [63:0] ap_return_49;
    output [63:0] ap_return_50;
    output [63:0] ap_return_51;
    output [63:0] ap_return_52;
    output [63:0] ap_return_53;
    output [63:0] ap_return_54;
    output [63:0] ap_return_55;
    output [63:0] ap_return_56;
    output [63:0] ap_return_57;
    output [63:0] ap_return_58;
    output [63:0] ap_return_59;
    output [63:0] ap_return_60;
    output [63:0] ap_return_61;
    output [63:0] ap_return_62;
    output [63:0] ap_return_63;

    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] p_read_17_reg_3029;
    reg   [63:0] p_read_17_reg_3029_pp0_iter1_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter2_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter3_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter4_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter5_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter6_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter7_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter8_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter9_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter10_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter11_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter12_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter13_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter14_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter15_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter16_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter17_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter18_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter19_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter20_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter21_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter22_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter23_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter24_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter25_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter26_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter27_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter28_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter29_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter30_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter31_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter32_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter33_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter34_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter35_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter36_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter37_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter38_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter39_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter40_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter41_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter42_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter43_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter44_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter45_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter46_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter47_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter48_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter49_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter50_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter51_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter52_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter53_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter54_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter55_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter56_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter57_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter58_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter59_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter60_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter61_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter62_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter63_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter64_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter65_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter66_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter67_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter68_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter69_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter70_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter71_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter72_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter73_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter74_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter75_reg;
    reg   [63:0] p_read_17_reg_3029_pp0_iter76_reg;
    reg   [63:0] p_read_18_reg_3034;
    reg   [63:0] p_read_18_reg_3034_pp0_iter1_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter2_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter3_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter4_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter5_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter6_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter7_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter8_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter9_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter10_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter11_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter12_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter13_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter14_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter15_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter16_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter17_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter18_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter19_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter20_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter21_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter22_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter23_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter24_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter25_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter26_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter27_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter28_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter29_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter30_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter31_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter32_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter33_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter34_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter35_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter36_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter37_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter38_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter39_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter40_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter41_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter42_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter43_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter44_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter45_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter46_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter47_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter48_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter49_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter50_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter51_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter52_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter53_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter54_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter55_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter56_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter57_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter58_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter59_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter60_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter61_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter62_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter63_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter64_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter65_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter66_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter67_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter68_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter69_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter70_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter71_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter72_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter73_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter74_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter75_reg;
    reg   [63:0] p_read_18_reg_3034_pp0_iter76_reg;
    reg   [63:0] p_read_19_reg_3039;
    reg   [63:0] p_read_19_reg_3039_pp0_iter1_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter2_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter3_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter4_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter5_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter6_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter7_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter8_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter9_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter10_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter11_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter12_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter13_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter14_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter15_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter16_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter17_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter18_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter19_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter20_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter21_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter22_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter23_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter24_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter25_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter26_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter27_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter28_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter29_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter30_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter31_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter32_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter33_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter34_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter35_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter36_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter37_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter38_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter39_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter40_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter41_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter42_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter43_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter44_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter45_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter46_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter47_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter48_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter49_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter50_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter51_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter52_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter53_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter54_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter55_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter56_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter57_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter58_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter59_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter60_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter61_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter62_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter63_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter64_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter65_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter66_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter67_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter68_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter69_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter70_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter71_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter72_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter73_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter74_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter75_reg;
    reg   [63:0] p_read_19_reg_3039_pp0_iter76_reg;
    reg   [63:0] p_read_20_reg_3044;
    reg   [63:0] p_read_20_reg_3044_pp0_iter1_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter2_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter3_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter4_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter5_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter6_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter7_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter8_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter9_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter10_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter11_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter12_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter13_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter14_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter15_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter16_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter17_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter18_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter19_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter20_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter21_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter22_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter23_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter24_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter25_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter26_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter27_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter28_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter29_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter30_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter31_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter32_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter33_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter34_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter35_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter36_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter37_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter38_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter39_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter40_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter41_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter42_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter43_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter44_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter45_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter46_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter47_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter48_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter49_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter50_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter51_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter52_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter53_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter54_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter55_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter56_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter57_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter58_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter59_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter60_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter61_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter62_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter63_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter64_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter65_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter66_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter67_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter68_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter69_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter70_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter71_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter72_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter73_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter74_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter75_reg;
    reg   [63:0] p_read_20_reg_3044_pp0_iter76_reg;
    reg   [63:0] p_read_21_reg_3049;
    reg   [63:0] p_read_21_reg_3049_pp0_iter1_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter2_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter3_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter4_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter5_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter6_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter7_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter8_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter9_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter10_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter11_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter12_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter13_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter14_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter15_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter16_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter17_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter18_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter19_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter20_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter21_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter22_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter23_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter24_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter25_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter26_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter27_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter28_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter29_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter30_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter31_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter32_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter33_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter34_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter35_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter36_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter37_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter38_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter39_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter40_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter41_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter42_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter43_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter44_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter45_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter46_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter47_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter48_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter49_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter50_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter51_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter52_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter53_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter54_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter55_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter56_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter57_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter58_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter59_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter60_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter61_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter62_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter63_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter64_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter65_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter66_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter67_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter68_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter69_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter70_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter71_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter72_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter73_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter74_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter75_reg;
    reg   [63:0] p_read_21_reg_3049_pp0_iter76_reg;
    reg   [63:0] p_read_22_reg_3054;
    reg   [63:0] p_read_22_reg_3054_pp0_iter1_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter2_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter3_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter4_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter5_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter6_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter7_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter8_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter9_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter10_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter11_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter12_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter13_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter14_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter15_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter16_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter17_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter18_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter19_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter20_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter21_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter22_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter23_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter24_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter25_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter26_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter27_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter28_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter29_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter30_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter31_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter32_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter33_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter34_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter35_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter36_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter37_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter38_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter39_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter40_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter41_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter42_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter43_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter44_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter45_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter46_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter47_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter48_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter49_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter50_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter51_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter52_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter53_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter54_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter55_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter56_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter57_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter58_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter59_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter60_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter61_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter62_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter63_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter64_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter65_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter66_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter67_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter68_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter69_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter70_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter71_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter72_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter73_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter74_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter75_reg;
    reg   [63:0] p_read_22_reg_3054_pp0_iter76_reg;
    reg   [63:0] p_read_23_reg_3059;
    reg   [63:0] p_read_23_reg_3059_pp0_iter1_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter2_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter3_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter4_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter5_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter6_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter7_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter8_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter9_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter10_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter11_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter12_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter13_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter14_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter15_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter16_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter17_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter18_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter19_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter20_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter21_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter22_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter23_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter24_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter25_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter26_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter27_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter28_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter29_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter30_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter31_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter32_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter33_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter34_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter35_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter36_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter37_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter38_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter39_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter40_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter41_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter42_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter43_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter44_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter45_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter46_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter47_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter48_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter49_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter50_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter51_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter52_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter53_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter54_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter55_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter56_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter57_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter58_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter59_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter60_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter61_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter62_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter63_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter64_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter65_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter66_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter67_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter68_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter69_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter70_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter71_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter72_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter73_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter74_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter75_reg;
    reg   [63:0] p_read_23_reg_3059_pp0_iter76_reg;
    reg   [63:0] p_read_24_reg_3064;
    reg   [63:0] p_read_24_reg_3064_pp0_iter1_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter2_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter3_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter4_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter5_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter6_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter7_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter8_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter9_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter10_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter11_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter12_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter13_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter14_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter15_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter16_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter17_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter18_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter19_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter20_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter21_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter22_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter23_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter24_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter25_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter26_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter27_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter28_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter29_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter30_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter31_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter32_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter33_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter34_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter35_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter36_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter37_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter38_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter39_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter40_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter41_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter42_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter43_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter44_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter45_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter46_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter47_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter48_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter49_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter50_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter51_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter52_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter53_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter54_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter55_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter56_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter57_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter58_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter59_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter60_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter61_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter62_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter63_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter64_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter65_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter66_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter67_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter68_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter69_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter70_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter71_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter72_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter73_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter74_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter75_reg;
    reg   [63:0] p_read_24_reg_3064_pp0_iter76_reg;
    reg   [63:0] p_read_25_reg_3069;
    reg   [63:0] p_read_25_reg_3069_pp0_iter1_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter2_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter3_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter4_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter5_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter6_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter7_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter8_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter9_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter10_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter11_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter12_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter13_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter14_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter15_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter16_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter17_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter18_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter19_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter20_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter21_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter22_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter23_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter24_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter25_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter26_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter27_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter28_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter29_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter30_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter31_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter32_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter33_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter34_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter35_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter36_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter37_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter38_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter39_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter40_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter41_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter42_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter43_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter44_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter45_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter46_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter47_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter48_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter49_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter50_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter51_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter52_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter53_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter54_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter55_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter56_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter57_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter58_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter59_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter60_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter61_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter62_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter63_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter64_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter65_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter66_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter67_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter68_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter69_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter70_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter71_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter72_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter73_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter74_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter75_reg;
    reg   [63:0] p_read_25_reg_3069_pp0_iter76_reg;
    reg   [63:0] p_read_26_reg_3074;
    reg   [63:0] p_read_26_reg_3074_pp0_iter1_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter2_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter3_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter4_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter5_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter6_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter7_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter8_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter9_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter10_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter11_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter12_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter13_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter14_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter15_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter16_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter17_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter18_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter19_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter20_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter21_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter22_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter23_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter24_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter25_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter26_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter27_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter28_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter29_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter30_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter31_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter32_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter33_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter34_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter35_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter36_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter37_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter38_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter39_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter40_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter41_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter42_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter43_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter44_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter45_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter46_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter47_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter48_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter49_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter50_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter51_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter52_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter53_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter54_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter55_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter56_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter57_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter58_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter59_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter60_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter61_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter62_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter63_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter64_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter65_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter66_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter67_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter68_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter69_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter70_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter71_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter72_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter73_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter74_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter75_reg;
    reg   [63:0] p_read_26_reg_3074_pp0_iter76_reg;
    reg   [63:0] p_read_27_reg_3079;
    reg   [63:0] p_read_27_reg_3079_pp0_iter1_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter2_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter3_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter4_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter5_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter6_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter7_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter8_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter9_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter10_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter11_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter12_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter13_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter14_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter15_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter16_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter17_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter18_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter19_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter20_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter21_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter22_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter23_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter24_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter25_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter26_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter27_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter28_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter29_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter30_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter31_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter32_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter33_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter34_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter35_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter36_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter37_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter38_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter39_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter40_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter41_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter42_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter43_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter44_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter45_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter46_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter47_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter48_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter49_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter50_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter51_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter52_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter53_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter54_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter55_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter56_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter57_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter58_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter59_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter60_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter61_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter62_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter63_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter64_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter65_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter66_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter67_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter68_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter69_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter70_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter71_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter72_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter73_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter74_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter75_reg;
    reg   [63:0] p_read_27_reg_3079_pp0_iter76_reg;
    reg   [63:0] p_read_28_reg_3084;
    reg   [63:0] p_read_28_reg_3084_pp0_iter1_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter2_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter3_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter4_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter5_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter6_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter7_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter8_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter9_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter10_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter11_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter12_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter13_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter14_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter15_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter16_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter17_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter18_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter19_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter20_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter21_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter22_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter23_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter24_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter25_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter26_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter27_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter28_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter29_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter30_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter31_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter32_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter33_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter34_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter35_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter36_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter37_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter38_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter39_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter40_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter41_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter42_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter43_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter44_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter45_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter46_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter47_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter48_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter49_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter50_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter51_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter52_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter53_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter54_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter55_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter56_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter57_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter58_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter59_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter60_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter61_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter62_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter63_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter64_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter65_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter66_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter67_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter68_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter69_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter70_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter71_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter72_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter73_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter74_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter75_reg;
    reg   [63:0] p_read_28_reg_3084_pp0_iter76_reg;
    reg   [63:0] p_read_29_reg_3089;
    reg   [63:0] p_read_29_reg_3089_pp0_iter1_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter2_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter3_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter4_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter5_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter6_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter7_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter8_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter9_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter10_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter11_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter12_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter13_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter14_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter15_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter16_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter17_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter18_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter19_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter20_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter21_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter22_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter23_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter24_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter25_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter26_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter27_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter28_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter29_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter30_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter31_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter32_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter33_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter34_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter35_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter36_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter37_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter38_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter39_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter40_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter41_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter42_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter43_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter44_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter45_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter46_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter47_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter48_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter49_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter50_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter51_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter52_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter53_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter54_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter55_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter56_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter57_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter58_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter59_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter60_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter61_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter62_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter63_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter64_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter65_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter66_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter67_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter68_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter69_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter70_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter71_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter72_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter73_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter74_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter75_reg;
    reg   [63:0] p_read_29_reg_3089_pp0_iter76_reg;
    reg   [63:0] p_read_30_reg_3094;
    reg   [63:0] p_read_30_reg_3094_pp0_iter1_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter2_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter3_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter4_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter5_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter6_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter7_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter8_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter9_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter10_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter11_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter12_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter13_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter14_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter15_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter16_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter17_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter18_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter19_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter20_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter21_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter22_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter23_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter24_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter25_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter26_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter27_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter28_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter29_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter30_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter31_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter32_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter33_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter34_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter35_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter36_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter37_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter38_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter39_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter40_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter41_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter42_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter43_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter44_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter45_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter46_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter47_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter48_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter49_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter50_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter51_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter52_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter53_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter54_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter55_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter56_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter57_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter58_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter59_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter60_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter61_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter62_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter63_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter64_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter65_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter66_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter67_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter68_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter69_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter70_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter71_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter72_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter73_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter74_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter75_reg;
    reg   [63:0] p_read_30_reg_3094_pp0_iter76_reg;
    reg   [63:0] p_read_31_reg_3099;
    reg   [63:0] p_read_31_reg_3099_pp0_iter1_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter2_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter3_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter4_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter5_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter6_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter7_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter8_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter9_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter10_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter11_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter12_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter13_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter14_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter15_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter16_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter17_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter18_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter19_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter20_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter21_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter22_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter23_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter24_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter25_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter26_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter27_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter28_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter29_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter30_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter31_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter32_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter33_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter34_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter35_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter36_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter37_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter38_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter39_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter40_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter41_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter42_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter43_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter44_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter45_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter46_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter47_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter48_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter49_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter50_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter51_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter52_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter53_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter54_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter55_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter56_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter57_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter58_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter59_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter60_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter61_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter62_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter63_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter64_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter65_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter66_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter67_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter68_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter69_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter70_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter71_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter72_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter73_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter74_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter75_reg;
    reg   [63:0] p_read_31_reg_3099_pp0_iter76_reg;
    reg   [63:0] p_read_32_reg_3104;
    reg   [63:0] p_read_32_reg_3104_pp0_iter1_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter2_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter3_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter4_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter5_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter6_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter7_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter8_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter9_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter10_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter11_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter12_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter13_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter14_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter15_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter16_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter17_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter18_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter19_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter20_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter21_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter22_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter23_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter24_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter25_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter26_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter27_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter28_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter29_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter30_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter31_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter32_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter33_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter34_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter35_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter36_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter37_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter38_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter39_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter40_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter41_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter42_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter43_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter44_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter45_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter46_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter47_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter48_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter49_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter50_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter51_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter52_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter53_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter54_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter55_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter56_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter57_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter58_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter59_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter60_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter61_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter62_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter63_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter64_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter65_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter66_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter67_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter68_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter69_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter70_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter71_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter72_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter73_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter74_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter75_reg;
    reg   [63:0] p_read_32_reg_3104_pp0_iter76_reg;
    reg   [63:0] p_read_33_reg_3109;
    reg   [63:0] p_read_33_reg_3109_pp0_iter1_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter2_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter3_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter4_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter5_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter6_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter7_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter8_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter9_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter10_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter11_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter12_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter13_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter14_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter15_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter16_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter17_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter18_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter19_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter20_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter21_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter22_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter23_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter24_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter25_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter26_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter27_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter28_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter29_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter30_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter31_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter32_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter33_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter34_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter35_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter36_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter37_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter38_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter39_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter40_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter41_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter42_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter43_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter44_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter45_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter46_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter47_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter48_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter49_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter50_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter51_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter52_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter53_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter54_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter55_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter56_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter57_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter58_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter59_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter60_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter61_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter62_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter63_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter64_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter65_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter66_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter67_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter68_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter69_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter70_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter71_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter72_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter73_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter74_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter75_reg;
    reg   [63:0] p_read_33_reg_3109_pp0_iter76_reg;
    reg   [63:0] p_read_34_reg_3114;
    reg   [63:0] p_read_34_reg_3114_pp0_iter1_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter2_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter3_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter4_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter5_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter6_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter7_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter8_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter9_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter10_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter11_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter12_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter13_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter14_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter15_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter16_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter17_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter18_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter19_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter20_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter21_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter22_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter23_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter24_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter25_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter26_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter27_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter28_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter29_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter30_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter31_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter32_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter33_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter34_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter35_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter36_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter37_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter38_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter39_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter40_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter41_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter42_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter43_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter44_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter45_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter46_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter47_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter48_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter49_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter50_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter51_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter52_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter53_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter54_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter55_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter56_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter57_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter58_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter59_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter60_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter61_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter62_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter63_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter64_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter65_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter66_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter67_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter68_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter69_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter70_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter71_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter72_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter73_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter74_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter75_reg;
    reg   [63:0] p_read_34_reg_3114_pp0_iter76_reg;
    reg   [63:0] p_read_35_reg_3119;
    reg   [63:0] p_read_35_reg_3119_pp0_iter1_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter2_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter3_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter4_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter5_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter6_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter7_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter8_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter9_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter10_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter11_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter12_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter13_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter14_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter15_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter16_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter17_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter18_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter19_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter20_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter21_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter22_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter23_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter24_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter25_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter26_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter27_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter28_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter29_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter30_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter31_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter32_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter33_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter34_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter35_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter36_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter37_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter38_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter39_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter40_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter41_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter42_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter43_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter44_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter45_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter46_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter47_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter48_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter49_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter50_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter51_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter52_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter53_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter54_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter55_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter56_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter57_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter58_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter59_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter60_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter61_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter62_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter63_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter64_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter65_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter66_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter67_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter68_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter69_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter70_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter71_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter72_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter73_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter74_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter75_reg;
    reg   [63:0] p_read_35_reg_3119_pp0_iter76_reg;
    reg   [63:0] p_read_36_reg_3124;
    reg   [63:0] p_read_36_reg_3124_pp0_iter1_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter2_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter3_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter4_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter5_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter6_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter7_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter8_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter9_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter10_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter11_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter12_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter13_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter14_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter15_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter16_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter17_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter18_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter19_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter20_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter21_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter22_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter23_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter24_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter25_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter26_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter27_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter28_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter29_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter30_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter31_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter32_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter33_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter34_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter35_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter36_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter37_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter38_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter39_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter40_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter41_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter42_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter43_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter44_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter45_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter46_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter47_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter48_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter49_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter50_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter51_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter52_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter53_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter54_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter55_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter56_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter57_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter58_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter59_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter60_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter61_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter62_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter63_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter64_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter65_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter66_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter67_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter68_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter69_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter70_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter71_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter72_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter73_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter74_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter75_reg;
    reg   [63:0] p_read_36_reg_3124_pp0_iter76_reg;
    reg   [63:0] p_read_37_reg_3129;
    reg   [63:0] p_read_37_reg_3129_pp0_iter1_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter2_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter3_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter4_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter5_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter6_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter7_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter8_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter9_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter10_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter11_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter12_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter13_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter14_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter15_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter16_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter17_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter18_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter19_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter20_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter21_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter22_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter23_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter24_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter25_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter26_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter27_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter28_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter29_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter30_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter31_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter32_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter33_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter34_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter35_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter36_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter37_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter38_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter39_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter40_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter41_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter42_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter43_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter44_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter45_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter46_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter47_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter48_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter49_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter50_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter51_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter52_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter53_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter54_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter55_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter56_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter57_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter58_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter59_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter60_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter61_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter62_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter63_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter64_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter65_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter66_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter67_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter68_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter69_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter70_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter71_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter72_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter73_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter74_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter75_reg;
    reg   [63:0] p_read_37_reg_3129_pp0_iter76_reg;
    reg   [63:0] p_read_38_reg_3134;
    reg   [63:0] p_read_38_reg_3134_pp0_iter1_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter2_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter3_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter4_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter5_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter6_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter7_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter8_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter9_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter10_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter11_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter12_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter13_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter14_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter15_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter16_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter17_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter18_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter19_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter20_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter21_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter22_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter23_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter24_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter25_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter26_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter27_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter28_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter29_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter30_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter31_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter32_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter33_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter34_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter35_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter36_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter37_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter38_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter39_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter40_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter41_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter42_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter43_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter44_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter45_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter46_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter47_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter48_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter49_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter50_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter51_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter52_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter53_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter54_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter55_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter56_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter57_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter58_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter59_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter60_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter61_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter62_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter63_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter64_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter65_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter66_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter67_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter68_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter69_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter70_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter71_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter72_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter73_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter74_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter75_reg;
    reg   [63:0] p_read_38_reg_3134_pp0_iter76_reg;
    reg   [63:0] p_read_39_reg_3139;
    reg   [63:0] p_read_39_reg_3139_pp0_iter1_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter2_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter3_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter4_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter5_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter6_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter7_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter8_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter9_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter10_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter11_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter12_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter13_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter14_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter15_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter16_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter17_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter18_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter19_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter20_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter21_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter22_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter23_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter24_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter25_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter26_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter27_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter28_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter29_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter30_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter31_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter32_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter33_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter34_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter35_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter36_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter37_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter38_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter39_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter40_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter41_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter42_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter43_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter44_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter45_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter46_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter47_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter48_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter49_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter50_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter51_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter52_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter53_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter54_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter55_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter56_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter57_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter58_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter59_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter60_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter61_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter62_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter63_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter64_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter65_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter66_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter67_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter68_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter69_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter70_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter71_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter72_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter73_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter74_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter75_reg;
    reg   [63:0] p_read_39_reg_3139_pp0_iter76_reg;
    reg   [63:0] p_read_40_reg_3144;
    reg   [63:0] p_read_40_reg_3144_pp0_iter1_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter2_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter3_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter4_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter5_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter6_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter7_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter8_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter9_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter10_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter11_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter12_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter13_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter14_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter15_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter16_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter17_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter18_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter19_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter20_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter21_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter22_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter23_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter24_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter25_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter26_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter27_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter28_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter29_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter30_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter31_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter32_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter33_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter34_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter35_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter36_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter37_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter38_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter39_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter40_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter41_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter42_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter43_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter44_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter45_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter46_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter47_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter48_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter49_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter50_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter51_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter52_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter53_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter54_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter55_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter56_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter57_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter58_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter59_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter60_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter61_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter62_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter63_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter64_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter65_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter66_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter67_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter68_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter69_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter70_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter71_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter72_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter73_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter74_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter75_reg;
    reg   [63:0] p_read_40_reg_3144_pp0_iter76_reg;
    reg   [63:0] p_read_41_reg_3149;
    reg   [63:0] p_read_41_reg_3149_pp0_iter1_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter2_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter3_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter4_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter5_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter6_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter7_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter8_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter9_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter10_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter11_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter12_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter13_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter14_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter15_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter16_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter17_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter18_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter19_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter20_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter21_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter22_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter23_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter24_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter25_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter26_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter27_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter28_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter29_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter30_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter31_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter32_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter33_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter34_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter35_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter36_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter37_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter38_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter39_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter40_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter41_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter42_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter43_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter44_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter45_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter46_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter47_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter48_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter49_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter50_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter51_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter52_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter53_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter54_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter55_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter56_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter57_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter58_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter59_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter60_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter61_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter62_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter63_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter64_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter65_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter66_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter67_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter68_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter69_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter70_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter71_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter72_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter73_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter74_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter75_reg;
    reg   [63:0] p_read_41_reg_3149_pp0_iter76_reg;
    reg   [63:0] p_read_42_reg_3154;
    reg   [63:0] p_read_42_reg_3154_pp0_iter1_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter2_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter3_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter4_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter5_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter6_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter7_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter8_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter9_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter10_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter11_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter12_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter13_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter14_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter15_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter16_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter17_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter18_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter19_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter20_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter21_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter22_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter23_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter24_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter25_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter26_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter27_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter28_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter29_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter30_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter31_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter32_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter33_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter34_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter35_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter36_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter37_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter38_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter39_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter40_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter41_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter42_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter43_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter44_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter45_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter46_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter47_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter48_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter49_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter50_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter51_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter52_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter53_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter54_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter55_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter56_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter57_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter58_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter59_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter60_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter61_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter62_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter63_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter64_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter65_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter66_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter67_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter68_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter69_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter70_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter71_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter72_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter73_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter74_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter75_reg;
    reg   [63:0] p_read_42_reg_3154_pp0_iter76_reg;
    reg   [63:0] p_read_43_reg_3159;
    reg   [63:0] p_read_43_reg_3159_pp0_iter1_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter2_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter3_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter4_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter5_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter6_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter7_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter8_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter9_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter10_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter11_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter12_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter13_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter14_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter15_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter16_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter17_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter18_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter19_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter20_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter21_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter22_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter23_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter24_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter25_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter26_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter27_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter28_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter29_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter30_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter31_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter32_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter33_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter34_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter35_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter36_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter37_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter38_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter39_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter40_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter41_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter42_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter43_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter44_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter45_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter46_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter47_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter48_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter49_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter50_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter51_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter52_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter53_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter54_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter55_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter56_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter57_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter58_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter59_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter60_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter61_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter62_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter63_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter64_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter65_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter66_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter67_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter68_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter69_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter70_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter71_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter72_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter73_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter74_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter75_reg;
    reg   [63:0] p_read_43_reg_3159_pp0_iter76_reg;
    reg   [63:0] p_read_44_reg_3164;
    reg   [63:0] p_read_44_reg_3164_pp0_iter1_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter2_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter3_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter4_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter5_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter6_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter7_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter8_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter9_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter10_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter11_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter12_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter13_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter14_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter15_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter16_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter17_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter18_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter19_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter20_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter21_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter22_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter23_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter24_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter25_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter26_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter27_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter28_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter29_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter30_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter31_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter32_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter33_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter34_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter35_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter36_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter37_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter38_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter39_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter40_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter41_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter42_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter43_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter44_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter45_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter46_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter47_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter48_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter49_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter50_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter51_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter52_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter53_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter54_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter55_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter56_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter57_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter58_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter59_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter60_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter61_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter62_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter63_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter64_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter65_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter66_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter67_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter68_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter69_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter70_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter71_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter72_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter73_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter74_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter75_reg;
    reg   [63:0] p_read_44_reg_3164_pp0_iter76_reg;
    reg   [63:0] p_read_45_reg_3169;
    reg   [63:0] p_read_45_reg_3169_pp0_iter1_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter2_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter3_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter4_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter5_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter6_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter7_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter8_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter9_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter10_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter11_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter12_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter13_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter14_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter15_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter16_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter17_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter18_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter19_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter20_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter21_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter22_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter23_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter24_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter25_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter26_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter27_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter28_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter29_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter30_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter31_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter32_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter33_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter34_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter35_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter36_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter37_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter38_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter39_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter40_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter41_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter42_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter43_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter44_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter45_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter46_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter47_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter48_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter49_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter50_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter51_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter52_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter53_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter54_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter55_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter56_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter57_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter58_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter59_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter60_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter61_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter62_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter63_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter64_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter65_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter66_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter67_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter68_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter69_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter70_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter71_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter72_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter73_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter74_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter75_reg;
    reg   [63:0] p_read_45_reg_3169_pp0_iter76_reg;
    reg   [63:0] p_read_46_reg_3174;
    reg   [63:0] p_read_46_reg_3174_pp0_iter1_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter2_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter3_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter4_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter5_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter6_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter7_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter8_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter9_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter10_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter11_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter12_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter13_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter14_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter15_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter16_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter17_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter18_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter19_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter20_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter21_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter22_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter23_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter24_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter25_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter26_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter27_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter28_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter29_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter30_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter31_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter32_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter33_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter34_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter35_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter36_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter37_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter38_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter39_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter40_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter41_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter42_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter43_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter44_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter45_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter46_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter47_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter48_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter49_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter50_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter51_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter52_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter53_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter54_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter55_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter56_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter57_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter58_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter59_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter60_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter61_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter62_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter63_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter64_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter65_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter66_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter67_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter68_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter69_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter70_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter71_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter72_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter73_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter74_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter75_reg;
    reg   [63:0] p_read_46_reg_3174_pp0_iter76_reg;
    reg   [63:0] p_read_47_reg_3179;
    reg   [63:0] p_read_47_reg_3179_pp0_iter1_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter2_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter3_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter4_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter5_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter6_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter7_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter8_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter9_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter10_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter11_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter12_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter13_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter14_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter15_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter16_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter17_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter18_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter19_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter20_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter21_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter22_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter23_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter24_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter25_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter26_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter27_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter28_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter29_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter30_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter31_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter32_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter33_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter34_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter35_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter36_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter37_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter38_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter39_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter40_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter41_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter42_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter43_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter44_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter45_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter46_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter47_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter48_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter49_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter50_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter51_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter52_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter53_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter54_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter55_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter56_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter57_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter58_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter59_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter60_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter61_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter62_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter63_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter64_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter65_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter66_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter67_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter68_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter69_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter70_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter71_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter72_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter73_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter74_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter75_reg;
    reg   [63:0] p_read_47_reg_3179_pp0_iter76_reg;
    reg   [63:0] p_read_48_reg_3184;
    reg   [63:0] p_read_48_reg_3184_pp0_iter1_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter2_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter3_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter4_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter5_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter6_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter7_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter8_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter9_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter10_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter11_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter12_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter13_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter14_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter15_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter16_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter17_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter18_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter19_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter20_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter21_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter22_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter23_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter24_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter25_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter26_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter27_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter28_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter29_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter30_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter31_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter32_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter33_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter34_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter35_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter36_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter37_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter38_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter39_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter40_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter41_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter42_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter43_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter44_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter45_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter46_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter47_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter48_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter49_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter50_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter51_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter52_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter53_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter54_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter55_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter56_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter57_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter58_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter59_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter60_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter61_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter62_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter63_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter64_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter65_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter66_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter67_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter68_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter69_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter70_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter71_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter72_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter73_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter74_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter75_reg;
    reg   [63:0] p_read_48_reg_3184_pp0_iter76_reg;
    reg   [63:0] p_read_49_reg_3189;
    reg   [63:0] p_read_49_reg_3189_pp0_iter1_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter2_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter3_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter4_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter5_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter6_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter7_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter8_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter9_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter10_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter11_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter12_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter13_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter14_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter15_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter16_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter17_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter18_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter19_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter20_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter21_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter22_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter23_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter24_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter25_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter26_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter27_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter28_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter29_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter30_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter31_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter32_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter33_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter34_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter35_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter36_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter37_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter38_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter39_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter40_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter41_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter42_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter43_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter44_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter45_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter46_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter47_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter48_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter49_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter50_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter51_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter52_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter53_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter54_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter55_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter56_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter57_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter58_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter59_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter60_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter61_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter62_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter63_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter64_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter65_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter66_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter67_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter68_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter69_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter70_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter71_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter72_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter73_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter74_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter75_reg;
    reg   [63:0] p_read_49_reg_3189_pp0_iter76_reg;
    reg   [63:0] p_read_50_reg_3194;
    reg   [63:0] p_read_50_reg_3194_pp0_iter1_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter2_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter3_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter4_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter5_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter6_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter7_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter8_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter9_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter10_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter11_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter12_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter13_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter14_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter15_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter16_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter17_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter18_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter19_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter20_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter21_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter22_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter23_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter24_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter25_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter26_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter27_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter28_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter29_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter30_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter31_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter32_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter33_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter34_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter35_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter36_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter37_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter38_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter39_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter40_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter41_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter42_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter43_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter44_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter45_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter46_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter47_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter48_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter49_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter50_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter51_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter52_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter53_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter54_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter55_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter56_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter57_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter58_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter59_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter60_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter61_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter62_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter63_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter64_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter65_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter66_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter67_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter68_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter69_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter70_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter71_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter72_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter73_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter74_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter75_reg;
    reg   [63:0] p_read_50_reg_3194_pp0_iter76_reg;
    reg   [63:0] p_read_51_reg_3199;
    reg   [63:0] p_read_51_reg_3199_pp0_iter1_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter2_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter3_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter4_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter5_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter6_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter7_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter8_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter9_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter10_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter11_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter12_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter13_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter14_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter15_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter16_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter17_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter18_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter19_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter20_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter21_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter22_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter23_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter24_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter25_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter26_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter27_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter28_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter29_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter30_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter31_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter32_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter33_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter34_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter35_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter36_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter37_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter38_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter39_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter40_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter41_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter42_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter43_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter44_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter45_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter46_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter47_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter48_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter49_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter50_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter51_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter52_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter53_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter54_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter55_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter56_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter57_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter58_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter59_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter60_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter61_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter62_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter63_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter64_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter65_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter66_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter67_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter68_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter69_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter70_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter71_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter72_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter73_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter74_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter75_reg;
    reg   [63:0] p_read_51_reg_3199_pp0_iter76_reg;
    reg   [63:0] p_read_52_reg_3204;
    reg   [63:0] p_read_52_reg_3204_pp0_iter1_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter2_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter3_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter4_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter5_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter6_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter7_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter8_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter9_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter10_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter11_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter12_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter13_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter14_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter15_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter16_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter17_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter18_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter19_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter20_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter21_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter22_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter23_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter24_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter25_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter26_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter27_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter28_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter29_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter30_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter31_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter32_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter33_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter34_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter35_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter36_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter37_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter38_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter39_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter40_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter41_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter42_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter43_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter44_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter45_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter46_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter47_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter48_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter49_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter50_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter51_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter52_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter53_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter54_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter55_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter56_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter57_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter58_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter59_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter60_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter61_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter62_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter63_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter64_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter65_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter66_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter67_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter68_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter69_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter70_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter71_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter72_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter73_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter74_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter75_reg;
    reg   [63:0] p_read_52_reg_3204_pp0_iter76_reg;
    reg   [63:0] p_read_53_reg_3209;
    reg   [63:0] p_read_53_reg_3209_pp0_iter1_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter2_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter3_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter4_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter5_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter6_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter7_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter8_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter9_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter10_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter11_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter12_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter13_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter14_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter15_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter16_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter17_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter18_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter19_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter20_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter21_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter22_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter23_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter24_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter25_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter26_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter27_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter28_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter29_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter30_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter31_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter32_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter33_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter34_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter35_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter36_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter37_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter38_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter39_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter40_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter41_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter42_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter43_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter44_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter45_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter46_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter47_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter48_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter49_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter50_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter51_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter52_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter53_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter54_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter55_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter56_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter57_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter58_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter59_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter60_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter61_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter62_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter63_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter64_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter65_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter66_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter67_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter68_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter69_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter70_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter71_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter72_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter73_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter74_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter75_reg;
    reg   [63:0] p_read_53_reg_3209_pp0_iter76_reg;
    reg   [63:0] p_read_54_reg_3214;
    reg   [63:0] p_read_54_reg_3214_pp0_iter1_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter2_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter3_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter4_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter5_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter6_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter7_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter8_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter9_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter10_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter11_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter12_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter13_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter14_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter15_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter16_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter17_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter18_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter19_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter20_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter21_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter22_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter23_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter24_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter25_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter26_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter27_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter28_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter29_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter30_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter31_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter32_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter33_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter34_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter35_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter36_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter37_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter38_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter39_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter40_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter41_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter42_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter43_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter44_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter45_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter46_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter47_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter48_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter49_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter50_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter51_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter52_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter53_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter54_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter55_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter56_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter57_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter58_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter59_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter60_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter61_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter62_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter63_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter64_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter65_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter66_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter67_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter68_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter69_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter70_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter71_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter72_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter73_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter74_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter75_reg;
    reg   [63:0] p_read_54_reg_3214_pp0_iter76_reg;
    reg   [63:0] p_read_55_reg_3219;
    reg   [63:0] p_read_55_reg_3219_pp0_iter1_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter2_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter3_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter4_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter5_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter6_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter7_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter8_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter9_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter10_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter11_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter12_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter13_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter14_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter15_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter16_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter17_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter18_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter19_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter20_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter21_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter22_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter23_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter24_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter25_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter26_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter27_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter28_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter29_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter30_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter31_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter32_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter33_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter34_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter35_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter36_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter37_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter38_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter39_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter40_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter41_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter42_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter43_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter44_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter45_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter46_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter47_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter48_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter49_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter50_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter51_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter52_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter53_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter54_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter55_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter56_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter57_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter58_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter59_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter60_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter61_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter62_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter63_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter64_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter65_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter66_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter67_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter68_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter69_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter70_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter71_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter72_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter73_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter74_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter75_reg;
    reg   [63:0] p_read_55_reg_3219_pp0_iter76_reg;
    reg   [63:0] p_read_56_reg_3224;
    reg   [63:0] p_read_56_reg_3224_pp0_iter1_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter2_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter3_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter4_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter5_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter6_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter7_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter8_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter9_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter10_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter11_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter12_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter13_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter14_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter15_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter16_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter17_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter18_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter19_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter20_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter21_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter22_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter23_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter24_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter25_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter26_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter27_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter28_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter29_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter30_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter31_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter32_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter33_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter34_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter35_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter36_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter37_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter38_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter39_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter40_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter41_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter42_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter43_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter44_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter45_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter46_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter47_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter48_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter49_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter50_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter51_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter52_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter53_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter54_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter55_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter56_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter57_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter58_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter59_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter60_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter61_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter62_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter63_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter64_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter65_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter66_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter67_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter68_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter69_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter70_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter71_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter72_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter73_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter74_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter75_reg;
    reg   [63:0] p_read_56_reg_3224_pp0_iter76_reg;
    reg   [63:0] p_read_57_reg_3229;
    reg   [63:0] p_read_57_reg_3229_pp0_iter1_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter2_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter3_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter4_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter5_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter6_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter7_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter8_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter9_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter10_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter11_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter12_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter13_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter14_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter15_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter16_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter17_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter18_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter19_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter20_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter21_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter22_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter23_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter24_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter25_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter26_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter27_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter28_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter29_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter30_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter31_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter32_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter33_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter34_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter35_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter36_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter37_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter38_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter39_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter40_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter41_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter42_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter43_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter44_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter45_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter46_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter47_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter48_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter49_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter50_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter51_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter52_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter53_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter54_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter55_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter56_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter57_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter58_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter59_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter60_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter61_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter62_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter63_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter64_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter65_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter66_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter67_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter68_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter69_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter70_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter71_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter72_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter73_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter74_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter75_reg;
    reg   [63:0] p_read_57_reg_3229_pp0_iter76_reg;
    reg   [63:0] p_read_58_reg_3234;
    reg   [63:0] p_read_58_reg_3234_pp0_iter1_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter2_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter3_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter4_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter5_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter6_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter7_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter8_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter9_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter10_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter11_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter12_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter13_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter14_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter15_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter16_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter17_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter18_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter19_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter20_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter21_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter22_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter23_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter24_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter25_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter26_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter27_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter28_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter29_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter30_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter31_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter32_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter33_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter34_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter35_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter36_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter37_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter38_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter39_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter40_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter41_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter42_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter43_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter44_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter45_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter46_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter47_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter48_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter49_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter50_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter51_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter52_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter53_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter54_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter55_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter56_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter57_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter58_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter59_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter60_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter61_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter62_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter63_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter64_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter65_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter66_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter67_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter68_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter69_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter70_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter71_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter72_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter73_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter74_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter75_reg;
    reg   [63:0] p_read_58_reg_3234_pp0_iter76_reg;
    reg   [63:0] p_read_59_reg_3239;
    reg   [63:0] p_read_59_reg_3239_pp0_iter1_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter2_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter3_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter4_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter5_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter6_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter7_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter8_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter9_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter10_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter11_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter12_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter13_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter14_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter15_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter16_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter17_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter18_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter19_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter20_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter21_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter22_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter23_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter24_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter25_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter26_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter27_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter28_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter29_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter30_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter31_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter32_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter33_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter34_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter35_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter36_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter37_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter38_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter39_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter40_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter41_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter42_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter43_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter44_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter45_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter46_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter47_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter48_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter49_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter50_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter51_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter52_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter53_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter54_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter55_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter56_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter57_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter58_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter59_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter60_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter61_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter62_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter63_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter64_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter65_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter66_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter67_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter68_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter69_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter70_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter71_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter72_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter73_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter74_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter75_reg;
    reg   [63:0] p_read_59_reg_3239_pp0_iter76_reg;
    reg   [63:0] p_read_60_reg_3244;
    reg   [63:0] p_read_60_reg_3244_pp0_iter1_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter2_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter3_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter4_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter5_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter6_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter7_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter8_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter9_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter10_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter11_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter12_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter13_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter14_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter15_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter16_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter17_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter18_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter19_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter20_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter21_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter22_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter23_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter24_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter25_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter26_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter27_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter28_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter29_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter30_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter31_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter32_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter33_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter34_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter35_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter36_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter37_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter38_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter39_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter40_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter41_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter42_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter43_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter44_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter45_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter46_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter47_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter48_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter49_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter50_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter51_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter52_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter53_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter54_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter55_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter56_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter57_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter58_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter59_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter60_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter61_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter62_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter63_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter64_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter65_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter66_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter67_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter68_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter69_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter70_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter71_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter72_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter73_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter74_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter75_reg;
    reg   [63:0] p_read_60_reg_3244_pp0_iter76_reg;
    reg   [63:0] p_read_61_reg_3249;
    reg   [63:0] p_read_61_reg_3249_pp0_iter1_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter2_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter3_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter4_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter5_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter6_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter7_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter8_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter9_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter10_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter11_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter12_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter13_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter14_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter15_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter16_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter17_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter18_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter19_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter20_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter21_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter22_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter23_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter24_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter25_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter26_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter27_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter28_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter29_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter30_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter31_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter32_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter33_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter34_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter35_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter36_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter37_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter38_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter39_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter40_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter41_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter42_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter43_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter44_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter45_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter46_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter47_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter48_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter49_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter50_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter51_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter52_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter53_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter54_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter55_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter56_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter57_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter58_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter59_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter60_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter61_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter62_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter63_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter64_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter65_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter66_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter67_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter68_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter69_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter70_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter71_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter72_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter73_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter74_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter75_reg;
    reg   [63:0] p_read_61_reg_3249_pp0_iter76_reg;
    reg   [63:0] p_read_62_reg_3254;
    reg   [63:0] p_read_62_reg_3254_pp0_iter1_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter2_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter3_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter4_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter5_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter6_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter7_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter8_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter9_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter10_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter11_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter12_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter13_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter14_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter15_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter16_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter17_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter18_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter19_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter20_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter21_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter22_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter23_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter24_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter25_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter26_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter27_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter28_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter29_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter30_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter31_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter32_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter33_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter34_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter35_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter36_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter37_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter38_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter39_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter40_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter41_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter42_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter43_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter44_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter45_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter46_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter47_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter48_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter49_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter50_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter51_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter52_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter53_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter54_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter55_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter56_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter57_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter58_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter59_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter60_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter61_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter62_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter63_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter64_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter65_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter66_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter67_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter68_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter69_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter70_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter71_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter72_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter73_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter74_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter75_reg;
    reg   [63:0] p_read_62_reg_3254_pp0_iter76_reg;
    reg   [63:0] p_read_63_reg_3259;
    reg   [63:0] p_read_63_reg_3259_pp0_iter1_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter2_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter3_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter4_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter5_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter6_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter7_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter8_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter9_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter10_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter11_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter12_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter13_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter14_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter15_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter16_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter17_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter18_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter19_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter20_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter21_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter22_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter23_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter24_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter25_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter26_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter27_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter28_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter29_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter30_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter31_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter32_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter33_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter34_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter35_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter36_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter37_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter38_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter39_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter40_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter41_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter42_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter43_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter44_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter45_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter46_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter47_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter48_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter49_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter50_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter51_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter52_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter53_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter54_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter55_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter56_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter57_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter58_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter59_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter60_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter61_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter62_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter63_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter64_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter65_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter66_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter67_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter68_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter69_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter70_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter71_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter72_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter73_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter74_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter75_reg;
    reg   [63:0] p_read_63_reg_3259_pp0_iter76_reg;
    reg   [63:0] p_read64_reg_3264;
    reg   [63:0] p_read64_reg_3264_pp0_iter1_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter2_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter3_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter4_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter5_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter6_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter7_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter8_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter9_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter10_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter11_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter12_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter13_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter14_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter15_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter16_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter17_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter18_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter19_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter20_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter21_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter22_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter23_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter24_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter25_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter26_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter27_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter28_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter29_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter30_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter31_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter32_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter33_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter34_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter35_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter36_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter37_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter38_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter39_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter40_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter41_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter42_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter43_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter44_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter45_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter46_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter47_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter48_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter49_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter50_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter51_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter52_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter53_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter54_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter55_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter56_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter57_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter58_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter59_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter60_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter61_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter62_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter63_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter64_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter65_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter66_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter67_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter68_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter69_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter70_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter71_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter72_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter73_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter74_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter75_reg;
    reg   [63:0] p_read64_reg_3264_pp0_iter76_reg;
    reg   [63:0] z_read_reg_3269;
    reg   [63:0] z_read_reg_3269_pp0_iter1_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter2_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter3_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter4_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter5_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter6_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter7_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter8_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter9_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter10_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter11_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter12_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter13_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter14_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter15_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter16_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter17_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter18_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter19_reg;
    reg   [63:0] z_read_reg_3269_pp0_iter20_reg;
    reg   [63:0] y_read_reg_3275;
    reg   [63:0] y_read_reg_3275_pp0_iter1_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter2_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter3_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter4_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter5_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter6_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter7_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter8_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter9_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter10_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter11_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter12_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter13_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter14_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter15_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter16_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter17_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter18_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter19_reg;
    reg   [63:0] y_read_reg_3275_pp0_iter20_reg;
    reg   [63:0] x_read_reg_3281;
    reg   [63:0] x_read_reg_3281_pp0_iter1_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter2_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter3_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter4_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter5_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter6_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter7_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter8_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter9_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter10_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter11_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter12_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter13_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter14_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter15_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter16_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter17_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter18_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter19_reg;
    reg   [63:0] x_read_reg_3281_pp0_iter20_reg;
    wire   [63:0] grp_fu_2089_p2;
    reg   [63:0] mul_i_0_0_3_reg_3287;
    wire   [63:0] grp_fu_2095_p2;
    reg   [63:0] mul_i_1_0_3_reg_3293;
    wire   [63:0] grp_fu_2101_p2;
    reg   [63:0] mul_i_2_0_3_reg_3299;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter7_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter8_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter9_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter10_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter11_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter12_reg;
    reg   [63:0] mul_i_2_0_3_reg_3299_pp0_iter13_reg;
    wire   [63:0] grp_fu_1718_p2;
    reg   [63:0] add_i_0_0_3_reg_3305;
    wire   [63:0] grp_fu_1723_p2;
    reg   [63:0] add_i_0_1_3_reg_3311;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter14_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter15_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter16_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter17_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter18_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter19_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter20_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter21_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter22_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter23_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter24_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter25_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter26_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter27_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter28_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter29_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter30_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter31_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter32_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter33_reg;
    reg   [63:0] add_i_0_1_3_reg_3311_pp0_iter34_reg;
    wire   [63:0] grp_fu_1728_p2;
    reg   [63:0] add_i_1_0_3_reg_3319;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter14_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter15_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter16_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter17_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter18_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter19_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter20_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter21_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter22_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter23_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter24_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter25_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter26_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter27_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter28_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter29_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter30_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter31_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter32_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter33_reg;
    reg   [63:0] add_i_1_0_3_reg_3319_pp0_iter34_reg;
    wire   [63:0] grp_fu_1733_p2;
    reg   [63:0] add_i_1_1_3_reg_3327;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter14_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter15_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter16_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter17_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter18_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter19_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter20_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter21_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter22_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter23_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter24_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter25_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter26_reg;
    reg   [63:0] add_i_1_1_3_reg_3327_pp0_iter27_reg;
    wire   [63:0] grp_fu_1738_p2;
    reg   [63:0] add_i_2_0_3_reg_3333;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter14_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter15_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter16_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter17_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter18_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter19_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter20_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter21_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter22_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter23_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter24_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter25_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter26_reg;
    reg   [63:0] add_i_2_0_3_reg_3333_pp0_iter27_reg;
    wire   [63:0] grp_fu_1743_p2;
    reg   [63:0] add_i_2_2_3_reg_3340;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter21_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter22_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter23_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter24_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter25_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter26_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter27_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter28_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter29_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter30_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter31_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter32_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter33_reg;
    reg   [63:0] add_i_2_2_3_reg_3340_pp0_iter34_reg;
    wire   [63:0] grp_fu_1748_p2;
    reg   [63:0] add_i1_reg_3347;
    wire   [63:0] grp_fu_2107_p2;
    reg   [63:0] mul_i1_0_0_1_reg_3352;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter21_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter22_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter23_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter24_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter25_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter26_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter27_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter28_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter29_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter30_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter31_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter32_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter33_reg;
    reg   [63:0] mul_i1_0_0_1_reg_3352_pp0_iter34_reg;
    wire   [63:0] grp_fu_2112_p2;
    reg   [63:0] mul_i1_0_1_reg_3360;
    wire   [63:0] grp_fu_2117_p2;
    reg   [63:0] mul_i1_1_0_1_reg_3365;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter21_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter22_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter23_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter24_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter25_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter26_reg;
    reg   [63:0] mul_i1_1_0_1_reg_3365_pp0_iter27_reg;
    wire   [63:0] grp_fu_2122_p2;
    reg   [63:0] mul_i1_1_1_reg_3371;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter21_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter22_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter23_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter24_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter25_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter26_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter27_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter28_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter29_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter30_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter31_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter32_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter33_reg;
    reg   [63:0] mul_i1_1_1_reg_3371_pp0_iter34_reg;
    wire   [63:0] grp_fu_2127_p2;
    reg   [63:0] mul_i1_2_0_1_reg_3378;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter21_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter22_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter23_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter24_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter25_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter26_reg;
    reg   [63:0] mul_i1_2_0_1_reg_3378_pp0_iter27_reg;
    wire   [63:0] grp_fu_1753_p2;
    reg   [63:0] add_i_0_3_3_reg_3385;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter28_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter29_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter30_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter31_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter32_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter33_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter34_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter35_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter36_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter37_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter38_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter39_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter40_reg;
    reg   [63:0] add_i_0_3_3_reg_3385_pp0_iter41_reg;
    wire   [63:0] grp_fu_1758_p2;
    reg   [63:0] add_i_1_3_3_reg_3391;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter28_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter29_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter30_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter31_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter32_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter33_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter34_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter35_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter36_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter37_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter38_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter39_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter40_reg;
    reg   [63:0] add_i_1_3_3_reg_3391_pp0_iter41_reg;
    wire   [63:0] grp_fu_1763_p2;
    reg   [63:0] add_i_2_3_3_reg_3397;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter28_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter29_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter30_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter31_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter32_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter33_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter34_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter35_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter36_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter37_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter38_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter39_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter40_reg;
    reg   [63:0] add_i_2_3_3_reg_3397_pp0_iter41_reg;
    wire   [63:0] grp_fu_1768_p2;
    reg   [63:0] add_i1_0_0_1_reg_3403;
    wire   [63:0] grp_fu_2132_p2;
    reg   [63:0] mul_i1_0_0_2_reg_3408;
    wire   [63:0] grp_fu_1772_p2;
    reg   [63:0] add_i1_0_1_reg_3413;
    wire   [63:0] grp_fu_1777_p2;
    reg   [63:0] add_i1_1_0_1_reg_3419;
    wire   [63:0] grp_fu_2137_p2;
    reg   [63:0] mul_i1_1_0_2_reg_3424;
    wire   [63:0] grp_fu_1781_p2;
    reg   [63:0] add_i1_1_1_reg_3429;
    wire   [63:0] grp_fu_1786_p2;
    reg   [63:0] add_i1_2_0_1_reg_3435;
    wire   [63:0] grp_fu_2142_p2;
    reg   [63:0] mul_i1_2_0_2_reg_3440;
    wire   [63:0] grp_fu_1790_p2;
    reg   [63:0] add_i1_2_1_reg_3445;
    wire   [63:0] grp_fu_1795_p2;
    reg   [63:0] add_i1_0_0_2_reg_3451;
    wire   [63:0] grp_fu_2147_p2;
    reg   [63:0] mul_i1_0_0_3_reg_3456;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter35_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter36_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter37_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter38_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter39_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter40_reg;
    reg   [63:0] mul_i1_0_0_3_reg_3456_pp0_iter41_reg;
    wire   [63:0] grp_fu_1799_p2;
    reg   [63:0] add_i1_0_1_1_reg_3463;
    wire   [63:0] grp_fu_1803_p2;
    reg   [63:0] add_i1_0_2_1_reg_3468;
    wire   [63:0] grp_fu_1807_p2;
    reg   [63:0] add_i1_1_0_2_reg_3474;
    wire   [63:0] grp_fu_2152_p2;
    reg   [63:0] mul_i1_1_0_3_reg_3479;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter35_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter36_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter37_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter38_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter39_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter40_reg;
    reg   [63:0] mul_i1_1_0_3_reg_3479_pp0_iter41_reg;
    wire   [63:0] grp_fu_1811_p2;
    reg   [63:0] add_i1_1_1_1_reg_3486;
    wire   [63:0] grp_fu_1815_p2;
    reg   [63:0] add_i1_1_2_1_reg_3491;
    wire   [63:0] grp_fu_1819_p2;
    reg   [63:0] add_i1_2_0_2_reg_3497;
    wire   [63:0] grp_fu_2157_p2;
    reg   [63:0] mul_i1_2_0_3_reg_3502;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter35_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter36_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter37_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter38_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter39_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter40_reg;
    reg   [63:0] mul_i1_2_0_3_reg_3502_pp0_iter41_reg;
    wire   [63:0] grp_fu_1823_p2;
    reg   [63:0] add_i1_2_1_1_reg_3509;
    wire   [63:0] grp_fu_2162_p2;
    reg   [63:0] mul_i1_2_1_2_reg_3514;
    wire   [63:0] grp_fu_1827_p2;
    reg   [63:0] add_i1_2_2_1_reg_3520;
    wire   [63:0] grp_fu_1831_p2;
    reg   [63:0] add_i1_0_0_3_reg_3526;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter42_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter43_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter44_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter45_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter46_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter47_reg;
    reg   [63:0] add_i1_0_0_3_reg_3526_pp0_iter48_reg;
    wire   [63:0] grp_fu_1835_p2;
    reg   [63:0] add_i1_0_1_2_reg_3532;
    wire   [63:0] grp_fu_1839_p2;
    reg   [63:0] add_i1_0_2_2_reg_3537;
    wire   [63:0] grp_fu_1843_p2;
    reg   [63:0] add_i1_0_3_2_reg_3542;
    wire   [63:0] grp_fu_1847_p2;
    reg   [63:0] add_i1_1_0_3_reg_3547;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter42_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter43_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter44_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter45_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter46_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter47_reg;
    reg   [63:0] add_i1_1_0_3_reg_3547_pp0_iter48_reg;
    wire   [63:0] grp_fu_1851_p2;
    reg   [63:0] add_i1_1_1_2_reg_3553;
    wire   [63:0] grp_fu_1855_p2;
    reg   [63:0] add_i1_1_2_2_reg_3558;
    wire   [63:0] grp_fu_1859_p2;
    reg   [63:0] add_i1_1_3_2_reg_3563;
    wire   [63:0] grp_fu_1863_p2;
    reg   [63:0] add_i1_2_0_3_reg_3568;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter42_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter43_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter44_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter45_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter46_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter47_reg;
    reg   [63:0] add_i1_2_0_3_reg_3568_pp0_iter48_reg;
    wire   [63:0] grp_fu_1867_p2;
    reg   [63:0] add_i1_2_1_2_reg_3574;
    wire   [63:0] grp_fu_1871_p2;
    reg   [63:0] add_i1_2_2_2_reg_3579;
    wire   [63:0] grp_fu_1875_p2;
    reg   [63:0] add_i1_2_3_2_reg_3584;
    wire   [63:0] grp_fu_1879_p2;
    reg   [63:0] add_i1_0_1_3_reg_3589;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter49_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter50_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter51_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter52_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter53_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter54_reg;
    reg   [63:0] add_i1_0_1_3_reg_3589_pp0_iter55_reg;
    wire   [63:0] grp_fu_1883_p2;
    reg   [63:0] add_i1_0_2_3_reg_3596;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter49_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter50_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter51_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter52_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter53_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter54_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter55_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter56_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter57_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter58_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter59_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter60_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter61_reg;
    reg   [63:0] add_i1_0_2_3_reg_3596_pp0_iter62_reg;
    wire   [63:0] grp_fu_1887_p2;
    reg   [63:0] add_i1_0_3_3_reg_3602;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter49_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter50_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter51_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter52_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter53_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter54_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter55_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter56_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter57_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter58_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter59_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter60_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter61_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter62_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter63_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter64_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter65_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter66_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter67_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter68_reg;
    reg   [63:0] add_i1_0_3_3_reg_3602_pp0_iter69_reg;
    wire   [63:0] grp_fu_1891_p2;
    reg   [63:0] add_i1_1_1_3_reg_3608;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter49_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter50_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter51_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter52_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter53_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter54_reg;
    reg   [63:0] add_i1_1_1_3_reg_3608_pp0_iter55_reg;
    wire   [63:0] grp_fu_1895_p2;
    reg   [63:0] add_i1_1_2_3_reg_3615;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter49_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter50_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter51_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter52_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter53_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter54_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter55_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter56_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter57_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter58_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter59_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter60_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter61_reg;
    reg   [63:0] add_i1_1_2_3_reg_3615_pp0_iter62_reg;
    wire   [63:0] grp_fu_1899_p2;
    reg   [63:0] add_i1_1_3_3_reg_3621;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter49_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter50_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter51_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter52_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter53_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter54_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter55_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter56_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter57_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter58_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter59_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter60_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter61_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter62_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter63_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter64_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter65_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter66_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter67_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter68_reg;
    reg   [63:0] add_i1_1_3_3_reg_3621_pp0_iter69_reg;
    wire   [63:0] grp_fu_1903_p2;
    reg   [63:0] add_i1_2_1_3_reg_3627;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter49_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter50_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter51_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter52_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter53_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter54_reg;
    reg   [63:0] add_i1_2_1_3_reg_3627_pp0_iter55_reg;
    wire   [63:0] grp_fu_1907_p2;
    reg   [63:0] add_i1_2_2_3_reg_3634;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter49_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter50_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter51_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter52_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter53_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter54_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter55_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter56_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter57_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter58_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter59_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter60_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter61_reg;
    reg   [63:0] add_i1_2_2_3_reg_3634_pp0_iter62_reg;
    wire   [63:0] grp_fu_1911_p2;
    reg   [63:0] add_i1_2_3_3_reg_3640;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter49_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter50_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter51_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter52_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter53_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter54_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter55_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter56_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter57_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter58_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter59_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter60_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter61_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter62_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter63_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter64_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter65_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter66_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter67_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter68_reg;
    reg   [63:0] add_i1_2_3_3_reg_3640_pp0_iter69_reg;
    wire   [63:0] grp_fu_2167_p2;
    reg   [63:0] mul_i2_0_1_reg_3646;
    wire   [63:0] grp_fu_2172_p2;
    reg   [63:0] mul_i2_1_1_reg_3651;
    wire   [63:0] grp_fu_2177_p2;
    reg   [63:0] mul_i2_2_1_reg_3656;
    wire   [63:0] grp_fu_1915_p2;
    reg   [63:0] add_i2_reg_3661;
    wire   [63:0] grp_fu_2182_p2;
    reg   [63:0] mul_i2_0_0_1_reg_3666;
    wire   [63:0] grp_fu_1920_p2;
    reg   [63:0] add_i2_0_1_reg_3672;
    wire   [63:0] grp_fu_2187_p2;
    reg   [63:0] mul_i2_0_2_1_reg_3679;
    wire   [63:0] grp_fu_1925_p2;
    reg   [63:0] add_i2_1_reg_3684;
    wire   [63:0] grp_fu_2192_p2;
    reg   [63:0] mul_i2_1_0_1_reg_3689;
    wire   [63:0] grp_fu_1930_p2;
    reg   [63:0] add_i2_1_1_reg_3695;
    wire   [63:0] grp_fu_2197_p2;
    reg   [63:0] mul_i2_1_2_1_reg_3702;
    wire   [63:0] grp_fu_1935_p2;
    reg   [63:0] add_i2_2_reg_3707;
    wire   [63:0] grp_fu_2202_p2;
    reg   [63:0] mul_i2_2_0_1_reg_3712;
    wire   [63:0] grp_fu_1940_p2;
    reg   [63:0] add_i2_2_1_reg_3718;
    wire   [63:0] grp_fu_2207_p2;
    reg   [63:0] mul_i2_2_2_1_reg_3725;
    wire   [63:0] grp_fu_1945_p2;
    reg   [63:0] add_i2_0_0_1_reg_3730;
    wire   [63:0] grp_fu_2212_p2;
    reg   [63:0] mul_i2_0_0_2_reg_3735;
    wire   [63:0] grp_fu_1949_p2;
    reg   [63:0] add_i2_0_1_1_reg_3742;
    wire   [63:0] grp_fu_1953_p2;
    reg   [63:0] add_i2_0_2_1_reg_3747;
    wire   [63:0] grp_fu_1957_p2;
    reg   [63:0] add_i2_0_3_1_reg_3752;
    wire   [63:0] grp_fu_1961_p2;
    reg   [63:0] add_i2_1_0_1_reg_3757;
    wire   [63:0] grp_fu_2217_p2;
    reg   [63:0] mul_i2_1_0_2_reg_3762;
    wire   [63:0] grp_fu_1965_p2;
    reg   [63:0] add_i2_1_1_1_reg_3769;
    wire   [63:0] grp_fu_1969_p2;
    reg   [63:0] add_i2_1_2_1_reg_3774;
    wire   [63:0] grp_fu_1973_p2;
    reg   [63:0] add_i2_1_3_1_reg_3779;
    wire   [63:0] grp_fu_1977_p2;
    reg   [63:0] add_i2_2_0_1_reg_3784;
    wire   [63:0] grp_fu_2222_p2;
    reg   [63:0] mul_i2_2_0_2_reg_3789;
    wire   [63:0] grp_fu_1981_p2;
    reg   [63:0] add_i2_2_1_1_reg_3796;
    wire   [63:0] grp_fu_1985_p2;
    reg   [63:0] add_i2_2_2_1_reg_3801;
    wire   [63:0] grp_fu_1989_p2;
    reg   [63:0] add_i2_2_3_1_reg_3806;
    wire   [63:0] grp_fu_1993_p2;
    reg   [63:0] add_i2_0_0_2_reg_3811;
    wire   [63:0] grp_fu_2227_p2;
    reg   [63:0] mul_i2_0_0_3_reg_3816;
    wire   [63:0] grp_fu_1997_p2;
    reg   [63:0] add_i2_0_1_2_reg_3823;
    wire   [63:0] grp_fu_2001_p2;
    reg   [63:0] add_i2_0_2_2_reg_3828;
    wire   [63:0] grp_fu_2005_p2;
    reg   [63:0] add_i2_0_3_2_reg_3833;
    wire   [63:0] grp_fu_2009_p2;
    reg   [63:0] add_i2_1_0_2_reg_3838;
    wire   [63:0] grp_fu_2232_p2;
    reg   [63:0] mul_i2_1_0_3_reg_3843;
    wire   [63:0] grp_fu_2013_p2;
    reg   [63:0] add_i2_1_1_2_reg_3850;
    wire   [63:0] grp_fu_2017_p2;
    reg   [63:0] add_i2_1_2_2_reg_3855;
    wire   [63:0] grp_fu_2021_p2;
    reg   [63:0] add_i2_1_3_2_reg_3860;
    wire   [63:0] grp_fu_2025_p2;
    reg   [63:0] add_i2_2_0_2_reg_3865;
    wire   [63:0] grp_fu_2237_p2;
    reg   [63:0] mul_i2_2_0_3_reg_3870;
    wire   [63:0] grp_fu_2029_p2;
    reg   [63:0] add_i2_2_1_2_reg_3877;
    wire   [63:0] grp_fu_2033_p2;
    reg   [63:0] add_i2_2_2_2_reg_3882;
    wire   [63:0] grp_fu_2037_p2;
    reg   [63:0] add_i2_2_3_2_reg_3887;
    wire   [63:0] grp_fu_2041_p2;
    reg   [63:0] H_0_03_reg_3892;
    wire   [63:0] grp_fu_2045_p2;
    reg   [63:0] H_0_16_reg_3900;
    wire   [63:0] grp_fu_2049_p2;
    reg   [63:0] H_0_27_reg_3908;
    wire   [63:0] grp_fu_2053_p2;
    reg   [63:0] H_0_3_reg_3916;
    wire   [63:0] grp_fu_2057_p2;
    reg   [63:0] H_1_0_reg_3924;
    wire   [63:0] grp_fu_2061_p2;
    reg   [63:0] H_1_1_reg_3932;
    wire   [63:0] grp_fu_2065_p2;
    reg   [63:0] H_1_2_reg_3940;
    wire   [63:0] grp_fu_2069_p2;
    reg   [63:0] H_1_3_reg_3948;
    wire   [63:0] grp_fu_2073_p2;
    reg   [63:0] H_2_0_reg_3956;
    wire   [63:0] grp_fu_2077_p2;
    reg   [63:0] H_2_1_reg_3964;
    wire   [63:0] grp_fu_2081_p2;
    reg   [63:0] H_2_2_reg_3972;
    wire   [63:0] grp_fu_2085_p2;
    reg   [63:0] H_2_3_reg_3980;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag11_0_reg_566;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag11_0_reg_566;
    wire   [1:0] H_offset_read_read_fu_158_p2;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag8_0_reg_585;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag8_0_reg_585;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag4_0_reg_604;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag4_0_reg_604;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag_0_reg_623;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag_0_reg_623;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag23_0_reg_642;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag23_0_reg_642;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag20_0_reg_661;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag20_0_reg_661;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag17_0_reg_680;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag17_0_reg_680;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag14_0_reg_699;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag14_0_reg_699;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag32_0_reg_718;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag32_0_reg_718;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag35_0_reg_737;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag35_0_reg_737;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag29_0_reg_756;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag29_0_reg_756;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag26_0_reg_775;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag26_0_reg_775;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag38_0_reg_794;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag38_0_reg_794;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag41_0_reg_813;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag41_0_reg_813;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag44_0_reg_832;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag44_0_reg_832;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag47_0_reg_851;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag47_0_reg_851;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag50_0_reg_870;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag50_0_reg_870;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag53_0_reg_889;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag53_0_reg_889;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag56_0_reg_908;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag56_0_reg_908;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag59_0_reg_927;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag59_0_reg_927;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag62_0_reg_946;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag62_0_reg_946;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag65_0_reg_965;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag65_0_reg_965;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag68_0_reg_984;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag68_0_reg_984;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag71_0_reg_1003;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag71_0_reg_1003;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag74_0_reg_1022;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag74_0_reg_1022;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag77_0_reg_1041;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag77_0_reg_1041;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag80_0_reg_1060;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag80_0_reg_1060;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag83_0_reg_1079;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag83_0_reg_1079;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag86_0_reg_1098;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag86_0_reg_1098;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag89_0_reg_1117;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag89_0_reg_1117;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag92_0_reg_1136;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag92_0_reg_1136;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag95_0_reg_1155;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag95_0_reg_1155;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag107_0_reg_1174;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag107_0_reg_1174;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag104_0_reg_1193;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag104_0_reg_1193;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag101_0_reg_1212;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag101_0_reg_1212;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag98_0_reg_1231;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag98_0_reg_1231;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag119_0_reg_1250;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag119_0_reg_1250;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag116_0_reg_1269;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag116_0_reg_1269;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag113_0_reg_1288;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag113_0_reg_1288;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag110_0_reg_1307;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag110_0_reg_1307;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag128_0_reg_1326;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag128_0_reg_1326;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag125_0_reg_1345;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag125_0_reg_1345;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag131_0_reg_1364;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag131_0_reg_1364;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag122_0_reg_1383;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag122_0_reg_1383;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag134_0_reg_1402;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag134_0_reg_1402;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag137_0_reg_1421;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag137_0_reg_1421;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag140_0_reg_1440;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag140_0_reg_1440;
    wire   [0:0] ap_phi_reg_pp0_iter0_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter1_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter2_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter3_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter4_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter5_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter6_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter7_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter8_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter9_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter10_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter11_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter12_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter13_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter14_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter15_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter16_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter17_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter18_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter19_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter20_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter21_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter22_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter23_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter24_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter25_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter26_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter27_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter28_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter29_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter30_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter31_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter32_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter33_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter34_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter35_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter36_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter37_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter38_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter39_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter40_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter41_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter42_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter43_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter44_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter45_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter46_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter47_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter48_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter49_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter50_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter51_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter52_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter53_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter54_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter55_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter56_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter57_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter58_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter59_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter60_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter61_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter62_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter63_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter64_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter65_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter66_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter67_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter68_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter69_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter70_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter71_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter72_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter73_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter74_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter75_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter76_write_flag143_0_reg_1459;
    reg   [0:0] ap_phi_reg_pp0_iter77_write_flag143_0_reg_1459;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_4_reg_1478;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_4_reg_1478;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_5_reg_1493;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_5_reg_1493;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_6_reg_1508;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_6_reg_1508;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_7_reg_1523;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_7_reg_1523;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_8_reg_1538;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_8_reg_1538;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_9_reg_1553;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_9_reg_1553;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_10_reg_1568;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_10_reg_1568;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_11_reg_1583;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_11_reg_1583;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_12_reg_1598;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_12_reg_1598;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_13_reg_1613;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_13_reg_1613;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_14_reg_1628;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_14_reg_1628;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_15_reg_1643;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_15_reg_1643;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_reg_1658;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_reg_1658;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_1_reg_1673;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_1_reg_1673;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_2_reg_1688;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_2_reg_1688;
    wire   [63:0] ap_phi_reg_pp0_iter0_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter1_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter2_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter3_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter4_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter5_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter6_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter7_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter8_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter9_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter10_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter11_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter12_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter13_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter14_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter15_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter16_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter17_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter18_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter19_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter20_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter21_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter22_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter23_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter24_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter25_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter26_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter27_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter28_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter29_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter30_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter31_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter32_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter33_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter34_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter35_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter36_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter37_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter38_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter39_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter40_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter41_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter42_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter43_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter44_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter45_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter46_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter47_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter48_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter49_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter50_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter51_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter52_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter53_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter54_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter55_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter56_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter57_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter58_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter59_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter60_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter61_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter62_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter63_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter64_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter65_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter66_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter67_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter68_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter69_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter70_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter71_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter72_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter73_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter74_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter75_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter76_phi_ln112_3_reg_1703;
    reg   [63:0] ap_phi_reg_pp0_iter77_phi_ln112_3_reg_1703;
    wire    ap_block_pp0_stage0;
    wire   [63:0] select_ln112_fu_2242_p3;
    wire   [63:0] select_ln112_1_fu_2248_p3;
    wire   [63:0] select_ln112_2_fu_2254_p3;
    wire   [63:0] select_ln112_3_fu_2260_p3;
    wire   [63:0] select_ln112_4_fu_2266_p3;
    wire   [63:0] select_ln112_5_fu_2272_p3;
    wire   [63:0] select_ln112_6_fu_2278_p3;
    wire   [63:0] select_ln112_7_fu_2284_p3;
    wire   [63:0] select_ln112_8_fu_2290_p3;
    wire   [63:0] select_ln112_9_fu_2296_p3;
    wire   [63:0] select_ln112_10_fu_2302_p3;
    wire   [63:0] select_ln112_11_fu_2308_p3;
    wire   [63:0] select_ln112_12_fu_2314_p3;
    wire   [63:0] select_ln112_13_fu_2320_p3;
    wire   [63:0] select_ln112_14_fu_2326_p3;
    wire   [63:0] select_ln112_15_fu_2332_p3;
    wire   [63:0] select_ln112_16_fu_2338_p3;
    wire   [63:0] select_ln112_17_fu_2344_p3;
    wire   [63:0] select_ln112_18_fu_2350_p3;
    wire   [63:0] select_ln112_19_fu_2356_p3;
    wire   [63:0] select_ln112_20_fu_2362_p3;
    wire   [63:0] select_ln112_21_fu_2368_p3;
    wire   [63:0] select_ln112_22_fu_2374_p3;
    wire   [63:0] select_ln112_23_fu_2380_p3;
    wire   [63:0] select_ln112_24_fu_2386_p3;
    wire   [63:0] select_ln112_25_fu_2392_p3;
    wire   [63:0] select_ln112_26_fu_2398_p3;
    wire   [63:0] select_ln112_27_fu_2404_p3;
    wire   [63:0] select_ln112_28_fu_2410_p3;
    wire   [63:0] select_ln112_29_fu_2416_p3;
    wire   [63:0] select_ln112_30_fu_2422_p3;
    wire   [63:0] select_ln112_31_fu_2428_p3;
    wire   [63:0] select_ln112_32_fu_2434_p3;
    wire   [63:0] select_ln112_33_fu_2440_p3;
    wire   [63:0] select_ln112_34_fu_2446_p3;
    wire   [63:0] select_ln112_35_fu_2452_p3;
    wire   [63:0] select_ln112_36_fu_2458_p3;
    wire   [63:0] select_ln112_37_fu_2464_p3;
    wire   [63:0] select_ln112_38_fu_2470_p3;
    wire   [63:0] select_ln112_39_fu_2476_p3;
    wire   [63:0] select_ln112_40_fu_2482_p3;
    wire   [63:0] select_ln112_41_fu_2488_p3;
    wire   [63:0] select_ln112_42_fu_2494_p3;
    wire   [63:0] select_ln112_43_fu_2500_p3;
    wire   [63:0] select_ln112_44_fu_2506_p3;
    wire   [63:0] select_ln112_45_fu_2512_p3;
    wire   [63:0] select_ln112_46_fu_2518_p3;
    wire   [63:0] select_ln112_47_fu_2524_p3;
    reg   [63:0] x_int_reg;
    reg   [63:0] y_int_reg;
    reg   [63:0] z_int_reg;
    reg   [63:0] p_read_int_reg;
    reg   [63:0] p_read1_int_reg;
    reg   [63:0] p_read2_int_reg;
    reg   [63:0] p_read3_int_reg;
    reg   [63:0] p_read4_int_reg;
    reg   [63:0] p_read5_int_reg;
    reg   [63:0] p_read6_int_reg;
    reg   [63:0] p_read7_int_reg;
    reg   [63:0] p_read8_int_reg;
    reg   [63:0] p_read9_int_reg;
    reg   [63:0] p_read10_int_reg;
    reg   [63:0] p_read11_int_reg;
    reg   [63:0] p_read12_int_reg;
    reg   [63:0] p_read13_int_reg;
    reg   [63:0] p_read14_int_reg;
    reg   [63:0] p_read15_int_reg;
    reg   [63:0] p_read16_int_reg;
    reg   [63:0] p_read17_int_reg;
    reg   [63:0] p_read18_int_reg;
    reg   [63:0] p_read19_int_reg;
    reg   [63:0] p_read20_int_reg;
    reg   [63:0] p_read21_int_reg;
    reg   [63:0] p_read22_int_reg;
    reg   [63:0] p_read23_int_reg;
    reg   [63:0] p_read24_int_reg;
    reg   [63:0] p_read25_int_reg;
    reg   [63:0] p_read26_int_reg;
    reg   [63:0] p_read27_int_reg;
    reg   [63:0] p_read28_int_reg;
    reg   [63:0] p_read29_int_reg;
    reg   [63:0] p_read30_int_reg;
    reg   [63:0] p_read31_int_reg;
    reg   [63:0] p_read32_int_reg;
    reg   [63:0] p_read33_int_reg;
    reg   [63:0] p_read34_int_reg;
    reg   [63:0] p_read35_int_reg;
    reg   [63:0] p_read36_int_reg;
    reg   [63:0] p_read37_int_reg;
    reg   [63:0] p_read38_int_reg;
    reg   [63:0] p_read39_int_reg;
    reg   [63:0] p_read40_int_reg;
    reg   [63:0] p_read41_int_reg;
    reg   [63:0] p_read42_int_reg;
    reg   [63:0] p_read43_int_reg;
    reg   [63:0] p_read44_int_reg;
    reg   [63:0] p_read45_int_reg;
    reg   [63:0] p_read46_int_reg;
    reg   [63:0] p_read47_int_reg;
    reg   [63:0] p_read48_int_reg;
    reg   [63:0] p_read49_int_reg;
    reg   [63:0] p_read50_int_reg;
    reg   [63:0] p_read51_int_reg;
    reg   [63:0] p_read52_int_reg;
    reg   [63:0] p_read53_int_reg;
    reg   [63:0] p_read54_int_reg;
    reg   [63:0] p_read55_int_reg;
    reg   [63:0] p_read56_int_reg;
    reg   [63:0] p_read57_int_reg;
    reg   [63:0] p_read58_int_reg;
    reg   [63:0] p_read59_int_reg;
    reg   [63:0] p_read60_int_reg;
    reg   [63:0] p_read61_int_reg;
    reg   [63:0] p_read62_int_reg;
    reg   [63:0] p_read63_int_reg;
    reg   [1:0] H_offset_int_reg;
    wire    ap_ce_reg;

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U520 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_3287),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_1718_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U521 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_3287),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1723_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U522 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_1_0_3_reg_3293),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1728_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U523 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_1_0_3_reg_3293),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_1733_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U524 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_2_0_3_reg_3299),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1738_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U525 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_2_0_3_reg_3299_pp0_iter13_reg),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_1743_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U526 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_3305),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1748_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U527 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x_read_reg_3281_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1753_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U528 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(y_read_reg_3275_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1758_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U529 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(z_read_reg_3269_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1763_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U530 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_reg_3347),
        .din1(mul_i1_0_0_1_reg_3352),
        .ce(1'b1),
        .dout(grp_fu_1768_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U531 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_0_1_reg_3360),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1772_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U532 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_3319_pp0_iter20_reg),
        .din1(mul_i1_1_0_1_reg_3365),
        .ce(1'b1),
        .dout(grp_fu_1777_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U533 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_1_1_reg_3371),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1781_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U534 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_0_3_reg_3333_pp0_iter20_reg),
        .din1(mul_i1_2_0_1_reg_3378),
        .ce(1'b1),
        .dout(grp_fu_1786_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U535 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_2_0_1_reg_3378),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1790_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U536 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_1_reg_3403),
        .din1(mul_i1_0_0_2_reg_3408),
        .ce(1'b1),
        .dout(grp_fu_1795_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U537 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_3413),
        .din1(add_i_0_1_3_reg_3311_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1799_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U538 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_3413),
        .din1(mul_i1_0_0_1_reg_3352_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1803_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U539 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_1_reg_3419),
        .din1(mul_i1_1_0_2_reg_3424),
        .ce(1'b1),
        .dout(grp_fu_1807_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U540 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_3429),
        .din1(add_i_1_1_3_reg_3327_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1811_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U541 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_3429),
        .din1(mul_i1_1_0_1_reg_3365_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1815_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U542 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_1_reg_3435),
        .din1(mul_i1_2_0_2_reg_3440),
        .ce(1'b1),
        .dout(grp_fu_1819_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U543 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_reg_3445),
        .din1(add_i_2_0_3_reg_3333_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1823_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U544 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_reg_3445),
        .din1(mul_i1_2_0_1_reg_3378_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_1827_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U545 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_2_reg_3451),
        .din1(mul_i1_0_0_3_reg_3456),
        .ce(1'b1),
        .dout(grp_fu_1831_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U546 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_1_reg_3463),
        .din1(mul_i1_0_0_1_reg_3352_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1835_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U547 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_3468),
        .din1(add_i_0_1_3_reg_3311_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1839_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U548 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_3468),
        .din1(mul_i1_0_0_1_reg_3352_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1843_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U549 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_2_reg_3474),
        .din1(mul_i1_1_0_3_reg_3479),
        .ce(1'b1),
        .dout(grp_fu_1847_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U550 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_1_reg_3486),
        .din1(mul_i1_1_1_reg_3371_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1851_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U551 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_3491),
        .din1(add_i_1_0_3_reg_3319_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1855_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U552 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_3491),
        .din1(mul_i1_1_1_reg_3371_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1859_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U553 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_2_reg_3497),
        .din1(mul_i1_2_0_3_reg_3502),
        .ce(1'b1),
        .dout(grp_fu_1863_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U554 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_1_reg_3509),
        .din1(mul_i1_2_1_2_reg_3514),
        .ce(1'b1),
        .dout(grp_fu_1867_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U555 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_3520),
        .din1(add_i_2_2_3_reg_3340_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_1871_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U556 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_3520),
        .din1(mul_i1_2_1_2_reg_3514),
        .ce(1'b1),
        .dout(grp_fu_1875_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U557 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_2_reg_3532),
        .din1(mul_i1_0_0_3_reg_3456_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1879_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U558 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_2_reg_3537),
        .din1(mul_i1_0_0_3_reg_3456_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1883_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U559 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_2_reg_3542),
        .din1(add_i_0_3_3_reg_3385_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1887_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U560 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_2_reg_3553),
        .din1(mul_i1_1_0_3_reg_3479_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1891_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U561 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_2_reg_3558),
        .din1(mul_i1_1_0_3_reg_3479_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1895_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U562 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_2_reg_3563),
        .din1(add_i_1_3_3_reg_3391_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1899_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U563 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_2_reg_3574),
        .din1(mul_i1_2_0_3_reg_3502_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1903_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U564 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_2_reg_3579),
        .din1(mul_i1_2_0_3_reg_3502_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1907_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U565 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_2_reg_3584),
        .din1(add_i_2_3_3_reg_3397_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_1911_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U566 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_3526_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1915_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U567 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_0_1_reg_3646),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1920_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U568 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_3547_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1925_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U569 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_1_1_reg_3651),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1930_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U570 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_3568_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1935_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U571 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_2_1_reg_3656),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_1940_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U572 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_reg_3661),
        .din1(mul_i2_0_0_1_reg_3666),
        .ce(1'b1),
        .dout(grp_fu_1945_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U573 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_3672),
        .din1(add_i1_0_1_3_reg_3589_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_1949_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U574 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_3672),
        .din1(mul_i2_0_2_1_reg_3679),
        .ce(1'b1),
        .dout(grp_fu_1953_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U575 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_3672),
        .din1(mul_i2_0_0_1_reg_3666),
        .ce(1'b1),
        .dout(grp_fu_1957_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U576 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_reg_3684),
        .din1(mul_i2_1_0_1_reg_3689),
        .ce(1'b1),
        .dout(grp_fu_1961_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U577 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_3695),
        .din1(add_i1_1_1_3_reg_3608_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_1965_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U578 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_3695),
        .din1(mul_i2_1_2_1_reg_3702),
        .ce(1'b1),
        .dout(grp_fu_1969_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U579 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_3695),
        .din1(mul_i2_1_0_1_reg_3689),
        .ce(1'b1),
        .dout(grp_fu_1973_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U580 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_reg_3707),
        .din1(mul_i2_2_0_1_reg_3712),
        .ce(1'b1),
        .dout(grp_fu_1977_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U581 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_3718),
        .din1(add_i1_2_1_3_reg_3627_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_1981_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U582 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_3718),
        .din1(mul_i2_2_2_1_reg_3725),
        .ce(1'b1),
        .dout(grp_fu_1985_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U583 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_3718),
        .din1(mul_i2_2_0_1_reg_3712),
        .ce(1'b1),
        .dout(grp_fu_1989_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U584 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_1_reg_3730),
        .din1(mul_i2_0_0_2_reg_3735),
        .ce(1'b1),
        .dout(grp_fu_1993_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U585 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_1_reg_3742),
        .din1(mul_i2_0_0_2_reg_3735),
        .ce(1'b1),
        .dout(grp_fu_1997_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U586 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_1_reg_3747),
        .din1(add_i1_0_2_3_reg_3596_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_2001_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U587 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_1_reg_3752),
        .din1(mul_i2_0_0_2_reg_3735),
        .ce(1'b1),
        .dout(grp_fu_2005_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U588 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_1_reg_3757),
        .din1(mul_i2_1_0_2_reg_3762),
        .ce(1'b1),
        .dout(grp_fu_2009_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U589 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_1_reg_3769),
        .din1(mul_i2_1_0_2_reg_3762),
        .ce(1'b1),
        .dout(grp_fu_2013_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U590 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_1_reg_3774),
        .din1(add_i1_1_2_3_reg_3615_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_2017_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U591 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_1_reg_3779),
        .din1(mul_i2_1_0_2_reg_3762),
        .ce(1'b1),
        .dout(grp_fu_2021_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U592 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_1_reg_3784),
        .din1(mul_i2_2_0_2_reg_3789),
        .ce(1'b1),
        .dout(grp_fu_2025_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U593 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_1_reg_3796),
        .din1(mul_i2_2_0_2_reg_3789),
        .ce(1'b1),
        .dout(grp_fu_2029_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U594 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_1_reg_3801),
        .din1(add_i1_2_2_3_reg_3634_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_2033_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U595 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_1_reg_3806),
        .din1(mul_i2_2_0_2_reg_3789),
        .ce(1'b1),
        .dout(grp_fu_2037_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U596 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_2_reg_3811),
        .din1(mul_i2_0_0_3_reg_3816),
        .ce(1'b1),
        .dout(grp_fu_2041_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U597 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_2_reg_3823),
        .din1(mul_i2_0_0_3_reg_3816),
        .ce(1'b1),
        .dout(grp_fu_2045_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U598 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_2_reg_3828),
        .din1(mul_i2_0_0_3_reg_3816),
        .ce(1'b1),
        .dout(grp_fu_2049_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U599 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_2_reg_3833),
        .din1(add_i1_0_3_3_reg_3602_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_2053_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U600 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_2_reg_3838),
        .din1(mul_i2_1_0_3_reg_3843),
        .ce(1'b1),
        .dout(grp_fu_2057_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U601 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_2_reg_3850),
        .din1(mul_i2_1_0_3_reg_3843),
        .ce(1'b1),
        .dout(grp_fu_2061_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U602 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_2_reg_3855),
        .din1(mul_i2_1_0_3_reg_3843),
        .ce(1'b1),
        .dout(grp_fu_2065_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U603 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_2_reg_3860),
        .din1(add_i1_1_3_3_reg_3621_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_2069_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U604 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_2_reg_3865),
        .din1(mul_i2_2_0_3_reg_3870),
        .ce(1'b1),
        .dout(grp_fu_2073_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U605 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_2_reg_3877),
        .din1(mul_i2_2_0_3_reg_3870),
        .ce(1'b1),
        .dout(grp_fu_2077_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U606 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_2_reg_3882),
        .din1(mul_i2_2_0_3_reg_3870),
        .ce(1'b1),
        .dout(grp_fu_2081_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U607 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_2_reg_3887),
        .din1(add_i1_2_3_3_reg_3640_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_2085_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U608 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x_int_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2089_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U609 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(y_int_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2095_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U610 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(z_int_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2101_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U611 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_3311),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2107_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U612 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_3305),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2112_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U613 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_1_3_reg_3327),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2117_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U614 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_3319),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2122_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U615 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_0_3_reg_3333),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2127_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U616 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_3311_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2132_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U617 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_3319_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2137_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U618 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_2_3_reg_3340),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2142_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U619 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_3_3_reg_3385),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2147_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U620 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_3_3_reg_3391),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2152_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U621 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_3_3_reg_3397),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2157_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U622 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_2_3_reg_3340_pp0_iter27_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2162_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U623 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_3526),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2167_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U624 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_3547),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2172_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U625 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_3568),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2177_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U626 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_3589),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2182_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U627 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_3589),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2187_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U628 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_3608),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2192_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U629 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_3608),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2197_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U630 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_3627),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2202_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U631 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_3627),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_2207_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U632 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_3_reg_3596_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2212_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U633 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_3_reg_3615_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2217_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U634 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_3_reg_3634_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2222_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U635 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_3_reg_3602_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2227_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U636 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_3_reg_3621_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2232_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U637 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_3_reg_3640_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_2237_p2)
    );

    always @(posedge ap_clk) begin
        H_offset_int_reg <= H_offset;
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_10_reg_1568 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_10_reg_1568 <= p_read54_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter0_phi_ln112_10_reg_1568;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_11_reg_1583 <= p_read55_int_reg;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_11_reg_1583 <= 64'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter0_phi_ln112_11_reg_1583;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_12_reg_1598 <= 64'd0;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_12_reg_1598 <= p_read56_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter0_phi_ln112_12_reg_1598;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_13_reg_1613 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_13_reg_1613 <= p_read57_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter0_phi_ln112_13_reg_1613;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_14_reg_1628 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_14_reg_1628 <= p_read58_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter0_phi_ln112_14_reg_1628;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_15_reg_1643 <= p_read59_int_reg;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_15_reg_1643 <= 64'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter0_phi_ln112_15_reg_1643;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_1_reg_1673 <= 64'd4607182418800017408;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_1_reg_1673 <= p_read61_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter0_phi_ln112_1_reg_1673;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_2_reg_1688 <= 64'd4607182418800017408;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_2_reg_1688 <= p_read62_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter0_phi_ln112_2_reg_1688;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_3_reg_1703 <= p_read63_int_reg;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_3_reg_1703 <= 64'd4607182418800017408;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter0_phi_ln112_3_reg_1703;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_4_reg_1478 <= 64'd0;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_4_reg_1478 <= p_read48_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter0_phi_ln112_4_reg_1478;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_5_reg_1493 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_5_reg_1493 <= p_read49_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter0_phi_ln112_5_reg_1493;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_6_reg_1508 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_6_reg_1508 <= p_read50_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter0_phi_ln112_6_reg_1508;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_7_reg_1523 <= p_read51_int_reg;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_7_reg_1523 <= 64'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter0_phi_ln112_7_reg_1523;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_8_reg_1538 <= 64'd0;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_8_reg_1538 <= p_read52_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter0_phi_ln112_8_reg_1538;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_9_reg_1553 <= 64'd0;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_9_reg_1553 <= p_read53_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter0_phi_ln112_9_reg_1553;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_reg_1658 <= 64'd4607182418800017408;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_phi_ln112_reg_1658 <= p_read60_int_reg;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter0_phi_ln112_reg_1658;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag101_0_reg_1212 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag101_0_reg_1212 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter0_write_flag101_0_reg_1212;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag104_0_reg_1193 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag104_0_reg_1193 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter0_write_flag104_0_reg_1193;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag107_0_reg_1174 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag107_0_reg_1174 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter0_write_flag107_0_reg_1174;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag110_0_reg_1307 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag110_0_reg_1307 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter0_write_flag110_0_reg_1307;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag113_0_reg_1288 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag113_0_reg_1288 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter0_write_flag113_0_reg_1288;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag116_0_reg_1269 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag116_0_reg_1269 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter0_write_flag116_0_reg_1269;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag119_0_reg_1250 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag119_0_reg_1250 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter0_write_flag119_0_reg_1250;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag11_0_reg_566 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag11_0_reg_566 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter0_write_flag11_0_reg_566;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag122_0_reg_1383 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag122_0_reg_1383 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter0_write_flag122_0_reg_1383;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag125_0_reg_1345 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag125_0_reg_1345 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter0_write_flag125_0_reg_1345;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag128_0_reg_1326 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag128_0_reg_1326 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter0_write_flag128_0_reg_1326;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag131_0_reg_1364 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag131_0_reg_1364 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter0_write_flag131_0_reg_1364;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag134_0_reg_1402 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag134_0_reg_1402 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter0_write_flag134_0_reg_1402;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag137_0_reg_1421 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag137_0_reg_1421 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter0_write_flag137_0_reg_1421;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag140_0_reg_1440 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag140_0_reg_1440 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter0_write_flag140_0_reg_1440;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag143_0_reg_1459 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag143_0_reg_1459 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter0_write_flag143_0_reg_1459;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag14_0_reg_699 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag14_0_reg_699 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter0_write_flag14_0_reg_699;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag17_0_reg_680 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag17_0_reg_680 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter0_write_flag17_0_reg_680;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag20_0_reg_661 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag20_0_reg_661 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter0_write_flag20_0_reg_661;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag23_0_reg_642 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag23_0_reg_642 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter0_write_flag23_0_reg_642;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag26_0_reg_775 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag26_0_reg_775 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter0_write_flag26_0_reg_775;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag29_0_reg_756 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag29_0_reg_756 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter0_write_flag29_0_reg_756;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag32_0_reg_718 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag32_0_reg_718 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter0_write_flag32_0_reg_718;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag35_0_reg_737 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag35_0_reg_737 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter0_write_flag35_0_reg_737;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag38_0_reg_794 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag38_0_reg_794 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter0_write_flag38_0_reg_794;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag41_0_reg_813 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag41_0_reg_813 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter0_write_flag41_0_reg_813;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag44_0_reg_832 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag44_0_reg_832 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter0_write_flag44_0_reg_832;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag47_0_reg_851 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag47_0_reg_851 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter0_write_flag47_0_reg_851;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag4_0_reg_604 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag4_0_reg_604 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter0_write_flag4_0_reg_604;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag50_0_reg_870 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag50_0_reg_870 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter0_write_flag50_0_reg_870;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag53_0_reg_889 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag53_0_reg_889 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter0_write_flag53_0_reg_889;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag56_0_reg_908 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag56_0_reg_908 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter0_write_flag56_0_reg_908;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag59_0_reg_927 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag59_0_reg_927 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter0_write_flag59_0_reg_927;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag62_0_reg_946 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag62_0_reg_946 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter0_write_flag62_0_reg_946;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag65_0_reg_965 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag65_0_reg_965 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter0_write_flag65_0_reg_965;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag68_0_reg_984 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag68_0_reg_984 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter0_write_flag68_0_reg_984;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag71_0_reg_1003 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag71_0_reg_1003 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter0_write_flag71_0_reg_1003;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag74_0_reg_1022 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag74_0_reg_1022 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter0_write_flag74_0_reg_1022;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag77_0_reg_1041 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag77_0_reg_1041 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter0_write_flag77_0_reg_1041;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag80_0_reg_1060 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag80_0_reg_1060 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter0_write_flag80_0_reg_1060;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag83_0_reg_1079 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag83_0_reg_1079 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter0_write_flag83_0_reg_1079;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag86_0_reg_1098 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag86_0_reg_1098 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter0_write_flag86_0_reg_1098;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag89_0_reg_1117 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag89_0_reg_1117 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter0_write_flag89_0_reg_1117;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag8_0_reg_585 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag8_0_reg_585 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter0_write_flag8_0_reg_585;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag92_0_reg_1136 <= 1'd1;
        end else if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag92_0_reg_1136 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter0_write_flag92_0_reg_1136;
        end
    end

    always @(posedge ap_clk) begin
        if ((((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag95_0_reg_1155 <= 1'd0;
        end else if (((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag95_0_reg_1155 <= 1'd1;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter0_write_flag95_0_reg_1155;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag98_0_reg_1231 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag98_0_reg_1231 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter0_write_flag98_0_reg_1231;
        end
    end

    always @(posedge ap_clk) begin
        if (((2'd0 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ap_phi_reg_pp0_iter1_write_flag_0_reg_623 <= 1'd1;
        end else if ((((2'd1 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd2 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)) | ((2'd3 == H_offset_read_read_fu_158_p2) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
            ap_phi_reg_pp0_iter1_write_flag_0_reg_623 <= 1'd0;
        end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            ap_phi_reg_pp0_iter1_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter0_write_flag_0_reg_623;
        end
    end

    always @(posedge ap_clk) begin
        p_read10_int_reg <= p_read10;
    end

    always @(posedge ap_clk) begin
        p_read11_int_reg <= p_read11;
    end

    always @(posedge ap_clk) begin
        p_read12_int_reg <= p_read12;
    end

    always @(posedge ap_clk) begin
        p_read13_int_reg <= p_read13;
    end

    always @(posedge ap_clk) begin
        p_read14_int_reg <= p_read14;
    end

    always @(posedge ap_clk) begin
        p_read15_int_reg <= p_read15;
    end

    always @(posedge ap_clk) begin
        p_read16_int_reg <= p_read16;
    end

    always @(posedge ap_clk) begin
        p_read17_int_reg <= p_read17;
    end

    always @(posedge ap_clk) begin
        p_read18_int_reg <= p_read18;
    end

    always @(posedge ap_clk) begin
        p_read19_int_reg <= p_read19;
    end

    always @(posedge ap_clk) begin
        p_read1_int_reg <= p_read1;
    end

    always @(posedge ap_clk) begin
        p_read20_int_reg <= p_read20;
    end

    always @(posedge ap_clk) begin
        p_read21_int_reg <= p_read21;
    end

    always @(posedge ap_clk) begin
        p_read22_int_reg <= p_read22;
    end

    always @(posedge ap_clk) begin
        p_read23_int_reg <= p_read23;
    end

    always @(posedge ap_clk) begin
        p_read24_int_reg <= p_read24;
    end

    always @(posedge ap_clk) begin
        p_read25_int_reg <= p_read25;
    end

    always @(posedge ap_clk) begin
        p_read26_int_reg <= p_read26;
    end

    always @(posedge ap_clk) begin
        p_read27_int_reg <= p_read27;
    end

    always @(posedge ap_clk) begin
        p_read28_int_reg <= p_read28;
    end

    always @(posedge ap_clk) begin
        p_read29_int_reg <= p_read29;
    end

    always @(posedge ap_clk) begin
        p_read2_int_reg <= p_read2;
    end

    always @(posedge ap_clk) begin
        p_read30_int_reg <= p_read30;
    end

    always @(posedge ap_clk) begin
        p_read31_int_reg <= p_read31;
    end

    always @(posedge ap_clk) begin
        p_read32_int_reg <= p_read32;
    end

    always @(posedge ap_clk) begin
        p_read33_int_reg <= p_read33;
    end

    always @(posedge ap_clk) begin
        p_read34_int_reg <= p_read34;
    end

    always @(posedge ap_clk) begin
        p_read35_int_reg <= p_read35;
    end

    always @(posedge ap_clk) begin
        p_read36_int_reg <= p_read36;
    end

    always @(posedge ap_clk) begin
        p_read37_int_reg <= p_read37;
    end

    always @(posedge ap_clk) begin
        p_read38_int_reg <= p_read38;
    end

    always @(posedge ap_clk) begin
        p_read39_int_reg <= p_read39;
    end

    always @(posedge ap_clk) begin
        p_read3_int_reg <= p_read3;
    end

    always @(posedge ap_clk) begin
        p_read40_int_reg <= p_read40;
    end

    always @(posedge ap_clk) begin
        p_read41_int_reg <= p_read41;
    end

    always @(posedge ap_clk) begin
        p_read42_int_reg <= p_read42;
    end

    always @(posedge ap_clk) begin
        p_read43_int_reg <= p_read43;
    end

    always @(posedge ap_clk) begin
        p_read44_int_reg <= p_read44;
    end

    always @(posedge ap_clk) begin
        p_read45_int_reg <= p_read45;
    end

    always @(posedge ap_clk) begin
        p_read46_int_reg <= p_read46;
    end

    always @(posedge ap_clk) begin
        p_read47_int_reg <= p_read47;
    end

    always @(posedge ap_clk) begin
        p_read48_int_reg <= p_read48;
    end

    always @(posedge ap_clk) begin
        p_read49_int_reg <= p_read49;
    end

    always @(posedge ap_clk) begin
        p_read4_int_reg <= p_read4;
    end

    always @(posedge ap_clk) begin
        p_read50_int_reg <= p_read50;
    end

    always @(posedge ap_clk) begin
        p_read51_int_reg <= p_read51;
    end

    always @(posedge ap_clk) begin
        p_read52_int_reg <= p_read52;
    end

    always @(posedge ap_clk) begin
        p_read53_int_reg <= p_read53;
    end

    always @(posedge ap_clk) begin
        p_read54_int_reg <= p_read54;
    end

    always @(posedge ap_clk) begin
        p_read55_int_reg <= p_read55;
    end

    always @(posedge ap_clk) begin
        p_read56_int_reg <= p_read56;
    end

    always @(posedge ap_clk) begin
        p_read57_int_reg <= p_read57;
    end

    always @(posedge ap_clk) begin
        p_read58_int_reg <= p_read58;
    end

    always @(posedge ap_clk) begin
        p_read59_int_reg <= p_read59;
    end

    always @(posedge ap_clk) begin
        p_read5_int_reg <= p_read5;
    end

    always @(posedge ap_clk) begin
        p_read60_int_reg <= p_read60;
    end

    always @(posedge ap_clk) begin
        p_read61_int_reg <= p_read61;
    end

    always @(posedge ap_clk) begin
        p_read62_int_reg <= p_read62;
    end

    always @(posedge ap_clk) begin
        p_read63_int_reg <= p_read63;
    end

    always @(posedge ap_clk) begin
        p_read6_int_reg <= p_read6;
    end

    always @(posedge ap_clk) begin
        p_read7_int_reg <= p_read7;
    end

    always @(posedge ap_clk) begin
        p_read8_int_reg <= p_read8;
    end

    always @(posedge ap_clk) begin
        p_read9_int_reg <= p_read9;
    end

    always @(posedge ap_clk) begin
        p_read_int_reg <= p_read;
    end

    always @(posedge ap_clk) begin
        x_int_reg <= x;
    end

    always @(posedge ap_clk) begin
        y_int_reg <= y;
    end

    always @(posedge ap_clk) begin
        z_int_reg <= z;
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            H_0_03_reg_3892 <= grp_fu_2041_p2;
            H_0_16_reg_3900 <= grp_fu_2045_p2;
            H_0_27_reg_3908 <= grp_fu_2049_p2;
            H_0_3_reg_3916 <= grp_fu_2053_p2;
            H_1_0_reg_3924 <= grp_fu_2057_p2;
            H_1_1_reg_3932 <= grp_fu_2061_p2;
            H_1_2_reg_3940 <= grp_fu_2065_p2;
            H_1_3_reg_3948 <= grp_fu_2069_p2;
            H_2_0_reg_3956 <= grp_fu_2073_p2;
            H_2_1_reg_3964 <= grp_fu_2077_p2;
            H_2_2_reg_3972 <= grp_fu_2081_p2;
            H_2_3_reg_3980 <= grp_fu_2085_p2;
            add_i1_0_0_1_reg_3403 <= grp_fu_1768_p2;
            add_i1_0_0_2_reg_3451 <= grp_fu_1795_p2;
            add_i1_0_0_3_reg_3526 <= grp_fu_1831_p2;
            add_i1_0_0_3_reg_3526_pp0_iter42_reg <= add_i1_0_0_3_reg_3526;
            add_i1_0_0_3_reg_3526_pp0_iter43_reg <= add_i1_0_0_3_reg_3526_pp0_iter42_reg;
            add_i1_0_0_3_reg_3526_pp0_iter44_reg <= add_i1_0_0_3_reg_3526_pp0_iter43_reg;
            add_i1_0_0_3_reg_3526_pp0_iter45_reg <= add_i1_0_0_3_reg_3526_pp0_iter44_reg;
            add_i1_0_0_3_reg_3526_pp0_iter46_reg <= add_i1_0_0_3_reg_3526_pp0_iter45_reg;
            add_i1_0_0_3_reg_3526_pp0_iter47_reg <= add_i1_0_0_3_reg_3526_pp0_iter46_reg;
            add_i1_0_0_3_reg_3526_pp0_iter48_reg <= add_i1_0_0_3_reg_3526_pp0_iter47_reg;
            add_i1_0_1_1_reg_3463 <= grp_fu_1799_p2;
            add_i1_0_1_2_reg_3532 <= grp_fu_1835_p2;
            add_i1_0_1_3_reg_3589 <= grp_fu_1879_p2;
            add_i1_0_1_3_reg_3589_pp0_iter49_reg <= add_i1_0_1_3_reg_3589;
            add_i1_0_1_3_reg_3589_pp0_iter50_reg <= add_i1_0_1_3_reg_3589_pp0_iter49_reg;
            add_i1_0_1_3_reg_3589_pp0_iter51_reg <= add_i1_0_1_3_reg_3589_pp0_iter50_reg;
            add_i1_0_1_3_reg_3589_pp0_iter52_reg <= add_i1_0_1_3_reg_3589_pp0_iter51_reg;
            add_i1_0_1_3_reg_3589_pp0_iter53_reg <= add_i1_0_1_3_reg_3589_pp0_iter52_reg;
            add_i1_0_1_3_reg_3589_pp0_iter54_reg <= add_i1_0_1_3_reg_3589_pp0_iter53_reg;
            add_i1_0_1_3_reg_3589_pp0_iter55_reg <= add_i1_0_1_3_reg_3589_pp0_iter54_reg;
            add_i1_0_1_reg_3413 <= grp_fu_1772_p2;
            add_i1_0_2_1_reg_3468 <= grp_fu_1803_p2;
            add_i1_0_2_2_reg_3537 <= grp_fu_1839_p2;
            add_i1_0_2_3_reg_3596 <= grp_fu_1883_p2;
            add_i1_0_2_3_reg_3596_pp0_iter49_reg <= add_i1_0_2_3_reg_3596;
            add_i1_0_2_3_reg_3596_pp0_iter50_reg <= add_i1_0_2_3_reg_3596_pp0_iter49_reg;
            add_i1_0_2_3_reg_3596_pp0_iter51_reg <= add_i1_0_2_3_reg_3596_pp0_iter50_reg;
            add_i1_0_2_3_reg_3596_pp0_iter52_reg <= add_i1_0_2_3_reg_3596_pp0_iter51_reg;
            add_i1_0_2_3_reg_3596_pp0_iter53_reg <= add_i1_0_2_3_reg_3596_pp0_iter52_reg;
            add_i1_0_2_3_reg_3596_pp0_iter54_reg <= add_i1_0_2_3_reg_3596_pp0_iter53_reg;
            add_i1_0_2_3_reg_3596_pp0_iter55_reg <= add_i1_0_2_3_reg_3596_pp0_iter54_reg;
            add_i1_0_2_3_reg_3596_pp0_iter56_reg <= add_i1_0_2_3_reg_3596_pp0_iter55_reg;
            add_i1_0_2_3_reg_3596_pp0_iter57_reg <= add_i1_0_2_3_reg_3596_pp0_iter56_reg;
            add_i1_0_2_3_reg_3596_pp0_iter58_reg <= add_i1_0_2_3_reg_3596_pp0_iter57_reg;
            add_i1_0_2_3_reg_3596_pp0_iter59_reg <= add_i1_0_2_3_reg_3596_pp0_iter58_reg;
            add_i1_0_2_3_reg_3596_pp0_iter60_reg <= add_i1_0_2_3_reg_3596_pp0_iter59_reg;
            add_i1_0_2_3_reg_3596_pp0_iter61_reg <= add_i1_0_2_3_reg_3596_pp0_iter60_reg;
            add_i1_0_2_3_reg_3596_pp0_iter62_reg <= add_i1_0_2_3_reg_3596_pp0_iter61_reg;
            add_i1_0_3_2_reg_3542 <= grp_fu_1843_p2;
            add_i1_0_3_3_reg_3602 <= grp_fu_1887_p2;
            add_i1_0_3_3_reg_3602_pp0_iter49_reg <= add_i1_0_3_3_reg_3602;
            add_i1_0_3_3_reg_3602_pp0_iter50_reg <= add_i1_0_3_3_reg_3602_pp0_iter49_reg;
            add_i1_0_3_3_reg_3602_pp0_iter51_reg <= add_i1_0_3_3_reg_3602_pp0_iter50_reg;
            add_i1_0_3_3_reg_3602_pp0_iter52_reg <= add_i1_0_3_3_reg_3602_pp0_iter51_reg;
            add_i1_0_3_3_reg_3602_pp0_iter53_reg <= add_i1_0_3_3_reg_3602_pp0_iter52_reg;
            add_i1_0_3_3_reg_3602_pp0_iter54_reg <= add_i1_0_3_3_reg_3602_pp0_iter53_reg;
            add_i1_0_3_3_reg_3602_pp0_iter55_reg <= add_i1_0_3_3_reg_3602_pp0_iter54_reg;
            add_i1_0_3_3_reg_3602_pp0_iter56_reg <= add_i1_0_3_3_reg_3602_pp0_iter55_reg;
            add_i1_0_3_3_reg_3602_pp0_iter57_reg <= add_i1_0_3_3_reg_3602_pp0_iter56_reg;
            add_i1_0_3_3_reg_3602_pp0_iter58_reg <= add_i1_0_3_3_reg_3602_pp0_iter57_reg;
            add_i1_0_3_3_reg_3602_pp0_iter59_reg <= add_i1_0_3_3_reg_3602_pp0_iter58_reg;
            add_i1_0_3_3_reg_3602_pp0_iter60_reg <= add_i1_0_3_3_reg_3602_pp0_iter59_reg;
            add_i1_0_3_3_reg_3602_pp0_iter61_reg <= add_i1_0_3_3_reg_3602_pp0_iter60_reg;
            add_i1_0_3_3_reg_3602_pp0_iter62_reg <= add_i1_0_3_3_reg_3602_pp0_iter61_reg;
            add_i1_0_3_3_reg_3602_pp0_iter63_reg <= add_i1_0_3_3_reg_3602_pp0_iter62_reg;
            add_i1_0_3_3_reg_3602_pp0_iter64_reg <= add_i1_0_3_3_reg_3602_pp0_iter63_reg;
            add_i1_0_3_3_reg_3602_pp0_iter65_reg <= add_i1_0_3_3_reg_3602_pp0_iter64_reg;
            add_i1_0_3_3_reg_3602_pp0_iter66_reg <= add_i1_0_3_3_reg_3602_pp0_iter65_reg;
            add_i1_0_3_3_reg_3602_pp0_iter67_reg <= add_i1_0_3_3_reg_3602_pp0_iter66_reg;
            add_i1_0_3_3_reg_3602_pp0_iter68_reg <= add_i1_0_3_3_reg_3602_pp0_iter67_reg;
            add_i1_0_3_3_reg_3602_pp0_iter69_reg <= add_i1_0_3_3_reg_3602_pp0_iter68_reg;
            add_i1_1_0_1_reg_3419 <= grp_fu_1777_p2;
            add_i1_1_0_2_reg_3474 <= grp_fu_1807_p2;
            add_i1_1_0_3_reg_3547 <= grp_fu_1847_p2;
            add_i1_1_0_3_reg_3547_pp0_iter42_reg <= add_i1_1_0_3_reg_3547;
            add_i1_1_0_3_reg_3547_pp0_iter43_reg <= add_i1_1_0_3_reg_3547_pp0_iter42_reg;
            add_i1_1_0_3_reg_3547_pp0_iter44_reg <= add_i1_1_0_3_reg_3547_pp0_iter43_reg;
            add_i1_1_0_3_reg_3547_pp0_iter45_reg <= add_i1_1_0_3_reg_3547_pp0_iter44_reg;
            add_i1_1_0_3_reg_3547_pp0_iter46_reg <= add_i1_1_0_3_reg_3547_pp0_iter45_reg;
            add_i1_1_0_3_reg_3547_pp0_iter47_reg <= add_i1_1_0_3_reg_3547_pp0_iter46_reg;
            add_i1_1_0_3_reg_3547_pp0_iter48_reg <= add_i1_1_0_3_reg_3547_pp0_iter47_reg;
            add_i1_1_1_1_reg_3486 <= grp_fu_1811_p2;
            add_i1_1_1_2_reg_3553 <= grp_fu_1851_p2;
            add_i1_1_1_3_reg_3608 <= grp_fu_1891_p2;
            add_i1_1_1_3_reg_3608_pp0_iter49_reg <= add_i1_1_1_3_reg_3608;
            add_i1_1_1_3_reg_3608_pp0_iter50_reg <= add_i1_1_1_3_reg_3608_pp0_iter49_reg;
            add_i1_1_1_3_reg_3608_pp0_iter51_reg <= add_i1_1_1_3_reg_3608_pp0_iter50_reg;
            add_i1_1_1_3_reg_3608_pp0_iter52_reg <= add_i1_1_1_3_reg_3608_pp0_iter51_reg;
            add_i1_1_1_3_reg_3608_pp0_iter53_reg <= add_i1_1_1_3_reg_3608_pp0_iter52_reg;
            add_i1_1_1_3_reg_3608_pp0_iter54_reg <= add_i1_1_1_3_reg_3608_pp0_iter53_reg;
            add_i1_1_1_3_reg_3608_pp0_iter55_reg <= add_i1_1_1_3_reg_3608_pp0_iter54_reg;
            add_i1_1_1_reg_3429 <= grp_fu_1781_p2;
            add_i1_1_2_1_reg_3491 <= grp_fu_1815_p2;
            add_i1_1_2_2_reg_3558 <= grp_fu_1855_p2;
            add_i1_1_2_3_reg_3615 <= grp_fu_1895_p2;
            add_i1_1_2_3_reg_3615_pp0_iter49_reg <= add_i1_1_2_3_reg_3615;
            add_i1_1_2_3_reg_3615_pp0_iter50_reg <= add_i1_1_2_3_reg_3615_pp0_iter49_reg;
            add_i1_1_2_3_reg_3615_pp0_iter51_reg <= add_i1_1_2_3_reg_3615_pp0_iter50_reg;
            add_i1_1_2_3_reg_3615_pp0_iter52_reg <= add_i1_1_2_3_reg_3615_pp0_iter51_reg;
            add_i1_1_2_3_reg_3615_pp0_iter53_reg <= add_i1_1_2_3_reg_3615_pp0_iter52_reg;
            add_i1_1_2_3_reg_3615_pp0_iter54_reg <= add_i1_1_2_3_reg_3615_pp0_iter53_reg;
            add_i1_1_2_3_reg_3615_pp0_iter55_reg <= add_i1_1_2_3_reg_3615_pp0_iter54_reg;
            add_i1_1_2_3_reg_3615_pp0_iter56_reg <= add_i1_1_2_3_reg_3615_pp0_iter55_reg;
            add_i1_1_2_3_reg_3615_pp0_iter57_reg <= add_i1_1_2_3_reg_3615_pp0_iter56_reg;
            add_i1_1_2_3_reg_3615_pp0_iter58_reg <= add_i1_1_2_3_reg_3615_pp0_iter57_reg;
            add_i1_1_2_3_reg_3615_pp0_iter59_reg <= add_i1_1_2_3_reg_3615_pp0_iter58_reg;
            add_i1_1_2_3_reg_3615_pp0_iter60_reg <= add_i1_1_2_3_reg_3615_pp0_iter59_reg;
            add_i1_1_2_3_reg_3615_pp0_iter61_reg <= add_i1_1_2_3_reg_3615_pp0_iter60_reg;
            add_i1_1_2_3_reg_3615_pp0_iter62_reg <= add_i1_1_2_3_reg_3615_pp0_iter61_reg;
            add_i1_1_3_2_reg_3563 <= grp_fu_1859_p2;
            add_i1_1_3_3_reg_3621 <= grp_fu_1899_p2;
            add_i1_1_3_3_reg_3621_pp0_iter49_reg <= add_i1_1_3_3_reg_3621;
            add_i1_1_3_3_reg_3621_pp0_iter50_reg <= add_i1_1_3_3_reg_3621_pp0_iter49_reg;
            add_i1_1_3_3_reg_3621_pp0_iter51_reg <= add_i1_1_3_3_reg_3621_pp0_iter50_reg;
            add_i1_1_3_3_reg_3621_pp0_iter52_reg <= add_i1_1_3_3_reg_3621_pp0_iter51_reg;
            add_i1_1_3_3_reg_3621_pp0_iter53_reg <= add_i1_1_3_3_reg_3621_pp0_iter52_reg;
            add_i1_1_3_3_reg_3621_pp0_iter54_reg <= add_i1_1_3_3_reg_3621_pp0_iter53_reg;
            add_i1_1_3_3_reg_3621_pp0_iter55_reg <= add_i1_1_3_3_reg_3621_pp0_iter54_reg;
            add_i1_1_3_3_reg_3621_pp0_iter56_reg <= add_i1_1_3_3_reg_3621_pp0_iter55_reg;
            add_i1_1_3_3_reg_3621_pp0_iter57_reg <= add_i1_1_3_3_reg_3621_pp0_iter56_reg;
            add_i1_1_3_3_reg_3621_pp0_iter58_reg <= add_i1_1_3_3_reg_3621_pp0_iter57_reg;
            add_i1_1_3_3_reg_3621_pp0_iter59_reg <= add_i1_1_3_3_reg_3621_pp0_iter58_reg;
            add_i1_1_3_3_reg_3621_pp0_iter60_reg <= add_i1_1_3_3_reg_3621_pp0_iter59_reg;
            add_i1_1_3_3_reg_3621_pp0_iter61_reg <= add_i1_1_3_3_reg_3621_pp0_iter60_reg;
            add_i1_1_3_3_reg_3621_pp0_iter62_reg <= add_i1_1_3_3_reg_3621_pp0_iter61_reg;
            add_i1_1_3_3_reg_3621_pp0_iter63_reg <= add_i1_1_3_3_reg_3621_pp0_iter62_reg;
            add_i1_1_3_3_reg_3621_pp0_iter64_reg <= add_i1_1_3_3_reg_3621_pp0_iter63_reg;
            add_i1_1_3_3_reg_3621_pp0_iter65_reg <= add_i1_1_3_3_reg_3621_pp0_iter64_reg;
            add_i1_1_3_3_reg_3621_pp0_iter66_reg <= add_i1_1_3_3_reg_3621_pp0_iter65_reg;
            add_i1_1_3_3_reg_3621_pp0_iter67_reg <= add_i1_1_3_3_reg_3621_pp0_iter66_reg;
            add_i1_1_3_3_reg_3621_pp0_iter68_reg <= add_i1_1_3_3_reg_3621_pp0_iter67_reg;
            add_i1_1_3_3_reg_3621_pp0_iter69_reg <= add_i1_1_3_3_reg_3621_pp0_iter68_reg;
            add_i1_2_0_1_reg_3435 <= grp_fu_1786_p2;
            add_i1_2_0_2_reg_3497 <= grp_fu_1819_p2;
            add_i1_2_0_3_reg_3568 <= grp_fu_1863_p2;
            add_i1_2_0_3_reg_3568_pp0_iter42_reg <= add_i1_2_0_3_reg_3568;
            add_i1_2_0_3_reg_3568_pp0_iter43_reg <= add_i1_2_0_3_reg_3568_pp0_iter42_reg;
            add_i1_2_0_3_reg_3568_pp0_iter44_reg <= add_i1_2_0_3_reg_3568_pp0_iter43_reg;
            add_i1_2_0_3_reg_3568_pp0_iter45_reg <= add_i1_2_0_3_reg_3568_pp0_iter44_reg;
            add_i1_2_0_3_reg_3568_pp0_iter46_reg <= add_i1_2_0_3_reg_3568_pp0_iter45_reg;
            add_i1_2_0_3_reg_3568_pp0_iter47_reg <= add_i1_2_0_3_reg_3568_pp0_iter46_reg;
            add_i1_2_0_3_reg_3568_pp0_iter48_reg <= add_i1_2_0_3_reg_3568_pp0_iter47_reg;
            add_i1_2_1_1_reg_3509 <= grp_fu_1823_p2;
            add_i1_2_1_2_reg_3574 <= grp_fu_1867_p2;
            add_i1_2_1_3_reg_3627 <= grp_fu_1903_p2;
            add_i1_2_1_3_reg_3627_pp0_iter49_reg <= add_i1_2_1_3_reg_3627;
            add_i1_2_1_3_reg_3627_pp0_iter50_reg <= add_i1_2_1_3_reg_3627_pp0_iter49_reg;
            add_i1_2_1_3_reg_3627_pp0_iter51_reg <= add_i1_2_1_3_reg_3627_pp0_iter50_reg;
            add_i1_2_1_3_reg_3627_pp0_iter52_reg <= add_i1_2_1_3_reg_3627_pp0_iter51_reg;
            add_i1_2_1_3_reg_3627_pp0_iter53_reg <= add_i1_2_1_3_reg_3627_pp0_iter52_reg;
            add_i1_2_1_3_reg_3627_pp0_iter54_reg <= add_i1_2_1_3_reg_3627_pp0_iter53_reg;
            add_i1_2_1_3_reg_3627_pp0_iter55_reg <= add_i1_2_1_3_reg_3627_pp0_iter54_reg;
            add_i1_2_1_reg_3445 <= grp_fu_1790_p2;
            add_i1_2_2_1_reg_3520 <= grp_fu_1827_p2;
            add_i1_2_2_2_reg_3579 <= grp_fu_1871_p2;
            add_i1_2_2_3_reg_3634 <= grp_fu_1907_p2;
            add_i1_2_2_3_reg_3634_pp0_iter49_reg <= add_i1_2_2_3_reg_3634;
            add_i1_2_2_3_reg_3634_pp0_iter50_reg <= add_i1_2_2_3_reg_3634_pp0_iter49_reg;
            add_i1_2_2_3_reg_3634_pp0_iter51_reg <= add_i1_2_2_3_reg_3634_pp0_iter50_reg;
            add_i1_2_2_3_reg_3634_pp0_iter52_reg <= add_i1_2_2_3_reg_3634_pp0_iter51_reg;
            add_i1_2_2_3_reg_3634_pp0_iter53_reg <= add_i1_2_2_3_reg_3634_pp0_iter52_reg;
            add_i1_2_2_3_reg_3634_pp0_iter54_reg <= add_i1_2_2_3_reg_3634_pp0_iter53_reg;
            add_i1_2_2_3_reg_3634_pp0_iter55_reg <= add_i1_2_2_3_reg_3634_pp0_iter54_reg;
            add_i1_2_2_3_reg_3634_pp0_iter56_reg <= add_i1_2_2_3_reg_3634_pp0_iter55_reg;
            add_i1_2_2_3_reg_3634_pp0_iter57_reg <= add_i1_2_2_3_reg_3634_pp0_iter56_reg;
            add_i1_2_2_3_reg_3634_pp0_iter58_reg <= add_i1_2_2_3_reg_3634_pp0_iter57_reg;
            add_i1_2_2_3_reg_3634_pp0_iter59_reg <= add_i1_2_2_3_reg_3634_pp0_iter58_reg;
            add_i1_2_2_3_reg_3634_pp0_iter60_reg <= add_i1_2_2_3_reg_3634_pp0_iter59_reg;
            add_i1_2_2_3_reg_3634_pp0_iter61_reg <= add_i1_2_2_3_reg_3634_pp0_iter60_reg;
            add_i1_2_2_3_reg_3634_pp0_iter62_reg <= add_i1_2_2_3_reg_3634_pp0_iter61_reg;
            add_i1_2_3_2_reg_3584 <= grp_fu_1875_p2;
            add_i1_2_3_3_reg_3640 <= grp_fu_1911_p2;
            add_i1_2_3_3_reg_3640_pp0_iter49_reg <= add_i1_2_3_3_reg_3640;
            add_i1_2_3_3_reg_3640_pp0_iter50_reg <= add_i1_2_3_3_reg_3640_pp0_iter49_reg;
            add_i1_2_3_3_reg_3640_pp0_iter51_reg <= add_i1_2_3_3_reg_3640_pp0_iter50_reg;
            add_i1_2_3_3_reg_3640_pp0_iter52_reg <= add_i1_2_3_3_reg_3640_pp0_iter51_reg;
            add_i1_2_3_3_reg_3640_pp0_iter53_reg <= add_i1_2_3_3_reg_3640_pp0_iter52_reg;
            add_i1_2_3_3_reg_3640_pp0_iter54_reg <= add_i1_2_3_3_reg_3640_pp0_iter53_reg;
            add_i1_2_3_3_reg_3640_pp0_iter55_reg <= add_i1_2_3_3_reg_3640_pp0_iter54_reg;
            add_i1_2_3_3_reg_3640_pp0_iter56_reg <= add_i1_2_3_3_reg_3640_pp0_iter55_reg;
            add_i1_2_3_3_reg_3640_pp0_iter57_reg <= add_i1_2_3_3_reg_3640_pp0_iter56_reg;
            add_i1_2_3_3_reg_3640_pp0_iter58_reg <= add_i1_2_3_3_reg_3640_pp0_iter57_reg;
            add_i1_2_3_3_reg_3640_pp0_iter59_reg <= add_i1_2_3_3_reg_3640_pp0_iter58_reg;
            add_i1_2_3_3_reg_3640_pp0_iter60_reg <= add_i1_2_3_3_reg_3640_pp0_iter59_reg;
            add_i1_2_3_3_reg_3640_pp0_iter61_reg <= add_i1_2_3_3_reg_3640_pp0_iter60_reg;
            add_i1_2_3_3_reg_3640_pp0_iter62_reg <= add_i1_2_3_3_reg_3640_pp0_iter61_reg;
            add_i1_2_3_3_reg_3640_pp0_iter63_reg <= add_i1_2_3_3_reg_3640_pp0_iter62_reg;
            add_i1_2_3_3_reg_3640_pp0_iter64_reg <= add_i1_2_3_3_reg_3640_pp0_iter63_reg;
            add_i1_2_3_3_reg_3640_pp0_iter65_reg <= add_i1_2_3_3_reg_3640_pp0_iter64_reg;
            add_i1_2_3_3_reg_3640_pp0_iter66_reg <= add_i1_2_3_3_reg_3640_pp0_iter65_reg;
            add_i1_2_3_3_reg_3640_pp0_iter67_reg <= add_i1_2_3_3_reg_3640_pp0_iter66_reg;
            add_i1_2_3_3_reg_3640_pp0_iter68_reg <= add_i1_2_3_3_reg_3640_pp0_iter67_reg;
            add_i1_2_3_3_reg_3640_pp0_iter69_reg <= add_i1_2_3_3_reg_3640_pp0_iter68_reg;
            add_i1_reg_3347 <= grp_fu_1748_p2;
            add_i2_0_0_1_reg_3730 <= grp_fu_1945_p2;
            add_i2_0_0_2_reg_3811 <= grp_fu_1993_p2;
            add_i2_0_1_1_reg_3742 <= grp_fu_1949_p2;
            add_i2_0_1_2_reg_3823 <= grp_fu_1997_p2;
            add_i2_0_1_reg_3672 <= grp_fu_1920_p2;
            add_i2_0_2_1_reg_3747 <= grp_fu_1953_p2;
            add_i2_0_2_2_reg_3828 <= grp_fu_2001_p2;
            add_i2_0_3_1_reg_3752 <= grp_fu_1957_p2;
            add_i2_0_3_2_reg_3833 <= grp_fu_2005_p2;
            add_i2_1_0_1_reg_3757 <= grp_fu_1961_p2;
            add_i2_1_0_2_reg_3838 <= grp_fu_2009_p2;
            add_i2_1_1_1_reg_3769 <= grp_fu_1965_p2;
            add_i2_1_1_2_reg_3850 <= grp_fu_2013_p2;
            add_i2_1_1_reg_3695 <= grp_fu_1930_p2;
            add_i2_1_2_1_reg_3774 <= grp_fu_1969_p2;
            add_i2_1_2_2_reg_3855 <= grp_fu_2017_p2;
            add_i2_1_3_1_reg_3779 <= grp_fu_1973_p2;
            add_i2_1_3_2_reg_3860 <= grp_fu_2021_p2;
            add_i2_1_reg_3684 <= grp_fu_1925_p2;
            add_i2_2_0_1_reg_3784 <= grp_fu_1977_p2;
            add_i2_2_0_2_reg_3865 <= grp_fu_2025_p2;
            add_i2_2_1_1_reg_3796 <= grp_fu_1981_p2;
            add_i2_2_1_2_reg_3877 <= grp_fu_2029_p2;
            add_i2_2_1_reg_3718 <= grp_fu_1940_p2;
            add_i2_2_2_1_reg_3801 <= grp_fu_1985_p2;
            add_i2_2_2_2_reg_3882 <= grp_fu_2033_p2;
            add_i2_2_3_1_reg_3806 <= grp_fu_1989_p2;
            add_i2_2_3_2_reg_3887 <= grp_fu_2037_p2;
            add_i2_2_reg_3707 <= grp_fu_1935_p2;
            add_i2_reg_3661 <= grp_fu_1915_p2;
            add_i_0_0_3_reg_3305 <= grp_fu_1718_p2;
            add_i_0_1_3_reg_3311 <= grp_fu_1723_p2;
            add_i_0_1_3_reg_3311_pp0_iter14_reg <= add_i_0_1_3_reg_3311;
            add_i_0_1_3_reg_3311_pp0_iter15_reg <= add_i_0_1_3_reg_3311_pp0_iter14_reg;
            add_i_0_1_3_reg_3311_pp0_iter16_reg <= add_i_0_1_3_reg_3311_pp0_iter15_reg;
            add_i_0_1_3_reg_3311_pp0_iter17_reg <= add_i_0_1_3_reg_3311_pp0_iter16_reg;
            add_i_0_1_3_reg_3311_pp0_iter18_reg <= add_i_0_1_3_reg_3311_pp0_iter17_reg;
            add_i_0_1_3_reg_3311_pp0_iter19_reg <= add_i_0_1_3_reg_3311_pp0_iter18_reg;
            add_i_0_1_3_reg_3311_pp0_iter20_reg <= add_i_0_1_3_reg_3311_pp0_iter19_reg;
            add_i_0_1_3_reg_3311_pp0_iter21_reg <= add_i_0_1_3_reg_3311_pp0_iter20_reg;
            add_i_0_1_3_reg_3311_pp0_iter22_reg <= add_i_0_1_3_reg_3311_pp0_iter21_reg;
            add_i_0_1_3_reg_3311_pp0_iter23_reg <= add_i_0_1_3_reg_3311_pp0_iter22_reg;
            add_i_0_1_3_reg_3311_pp0_iter24_reg <= add_i_0_1_3_reg_3311_pp0_iter23_reg;
            add_i_0_1_3_reg_3311_pp0_iter25_reg <= add_i_0_1_3_reg_3311_pp0_iter24_reg;
            add_i_0_1_3_reg_3311_pp0_iter26_reg <= add_i_0_1_3_reg_3311_pp0_iter25_reg;
            add_i_0_1_3_reg_3311_pp0_iter27_reg <= add_i_0_1_3_reg_3311_pp0_iter26_reg;
            add_i_0_1_3_reg_3311_pp0_iter28_reg <= add_i_0_1_3_reg_3311_pp0_iter27_reg;
            add_i_0_1_3_reg_3311_pp0_iter29_reg <= add_i_0_1_3_reg_3311_pp0_iter28_reg;
            add_i_0_1_3_reg_3311_pp0_iter30_reg <= add_i_0_1_3_reg_3311_pp0_iter29_reg;
            add_i_0_1_3_reg_3311_pp0_iter31_reg <= add_i_0_1_3_reg_3311_pp0_iter30_reg;
            add_i_0_1_3_reg_3311_pp0_iter32_reg <= add_i_0_1_3_reg_3311_pp0_iter31_reg;
            add_i_0_1_3_reg_3311_pp0_iter33_reg <= add_i_0_1_3_reg_3311_pp0_iter32_reg;
            add_i_0_1_3_reg_3311_pp0_iter34_reg <= add_i_0_1_3_reg_3311_pp0_iter33_reg;
            add_i_0_3_3_reg_3385 <= grp_fu_1753_p2;
            add_i_0_3_3_reg_3385_pp0_iter28_reg <= add_i_0_3_3_reg_3385;
            add_i_0_3_3_reg_3385_pp0_iter29_reg <= add_i_0_3_3_reg_3385_pp0_iter28_reg;
            add_i_0_3_3_reg_3385_pp0_iter30_reg <= add_i_0_3_3_reg_3385_pp0_iter29_reg;
            add_i_0_3_3_reg_3385_pp0_iter31_reg <= add_i_0_3_3_reg_3385_pp0_iter30_reg;
            add_i_0_3_3_reg_3385_pp0_iter32_reg <= add_i_0_3_3_reg_3385_pp0_iter31_reg;
            add_i_0_3_3_reg_3385_pp0_iter33_reg <= add_i_0_3_3_reg_3385_pp0_iter32_reg;
            add_i_0_3_3_reg_3385_pp0_iter34_reg <= add_i_0_3_3_reg_3385_pp0_iter33_reg;
            add_i_0_3_3_reg_3385_pp0_iter35_reg <= add_i_0_3_3_reg_3385_pp0_iter34_reg;
            add_i_0_3_3_reg_3385_pp0_iter36_reg <= add_i_0_3_3_reg_3385_pp0_iter35_reg;
            add_i_0_3_3_reg_3385_pp0_iter37_reg <= add_i_0_3_3_reg_3385_pp0_iter36_reg;
            add_i_0_3_3_reg_3385_pp0_iter38_reg <= add_i_0_3_3_reg_3385_pp0_iter37_reg;
            add_i_0_3_3_reg_3385_pp0_iter39_reg <= add_i_0_3_3_reg_3385_pp0_iter38_reg;
            add_i_0_3_3_reg_3385_pp0_iter40_reg <= add_i_0_3_3_reg_3385_pp0_iter39_reg;
            add_i_0_3_3_reg_3385_pp0_iter41_reg <= add_i_0_3_3_reg_3385_pp0_iter40_reg;
            add_i_1_0_3_reg_3319 <= grp_fu_1728_p2;
            add_i_1_0_3_reg_3319_pp0_iter14_reg <= add_i_1_0_3_reg_3319;
            add_i_1_0_3_reg_3319_pp0_iter15_reg <= add_i_1_0_3_reg_3319_pp0_iter14_reg;
            add_i_1_0_3_reg_3319_pp0_iter16_reg <= add_i_1_0_3_reg_3319_pp0_iter15_reg;
            add_i_1_0_3_reg_3319_pp0_iter17_reg <= add_i_1_0_3_reg_3319_pp0_iter16_reg;
            add_i_1_0_3_reg_3319_pp0_iter18_reg <= add_i_1_0_3_reg_3319_pp0_iter17_reg;
            add_i_1_0_3_reg_3319_pp0_iter19_reg <= add_i_1_0_3_reg_3319_pp0_iter18_reg;
            add_i_1_0_3_reg_3319_pp0_iter20_reg <= add_i_1_0_3_reg_3319_pp0_iter19_reg;
            add_i_1_0_3_reg_3319_pp0_iter21_reg <= add_i_1_0_3_reg_3319_pp0_iter20_reg;
            add_i_1_0_3_reg_3319_pp0_iter22_reg <= add_i_1_0_3_reg_3319_pp0_iter21_reg;
            add_i_1_0_3_reg_3319_pp0_iter23_reg <= add_i_1_0_3_reg_3319_pp0_iter22_reg;
            add_i_1_0_3_reg_3319_pp0_iter24_reg <= add_i_1_0_3_reg_3319_pp0_iter23_reg;
            add_i_1_0_3_reg_3319_pp0_iter25_reg <= add_i_1_0_3_reg_3319_pp0_iter24_reg;
            add_i_1_0_3_reg_3319_pp0_iter26_reg <= add_i_1_0_3_reg_3319_pp0_iter25_reg;
            add_i_1_0_3_reg_3319_pp0_iter27_reg <= add_i_1_0_3_reg_3319_pp0_iter26_reg;
            add_i_1_0_3_reg_3319_pp0_iter28_reg <= add_i_1_0_3_reg_3319_pp0_iter27_reg;
            add_i_1_0_3_reg_3319_pp0_iter29_reg <= add_i_1_0_3_reg_3319_pp0_iter28_reg;
            add_i_1_0_3_reg_3319_pp0_iter30_reg <= add_i_1_0_3_reg_3319_pp0_iter29_reg;
            add_i_1_0_3_reg_3319_pp0_iter31_reg <= add_i_1_0_3_reg_3319_pp0_iter30_reg;
            add_i_1_0_3_reg_3319_pp0_iter32_reg <= add_i_1_0_3_reg_3319_pp0_iter31_reg;
            add_i_1_0_3_reg_3319_pp0_iter33_reg <= add_i_1_0_3_reg_3319_pp0_iter32_reg;
            add_i_1_0_3_reg_3319_pp0_iter34_reg <= add_i_1_0_3_reg_3319_pp0_iter33_reg;
            add_i_1_1_3_reg_3327 <= grp_fu_1733_p2;
            add_i_1_1_3_reg_3327_pp0_iter14_reg <= add_i_1_1_3_reg_3327;
            add_i_1_1_3_reg_3327_pp0_iter15_reg <= add_i_1_1_3_reg_3327_pp0_iter14_reg;
            add_i_1_1_3_reg_3327_pp0_iter16_reg <= add_i_1_1_3_reg_3327_pp0_iter15_reg;
            add_i_1_1_3_reg_3327_pp0_iter17_reg <= add_i_1_1_3_reg_3327_pp0_iter16_reg;
            add_i_1_1_3_reg_3327_pp0_iter18_reg <= add_i_1_1_3_reg_3327_pp0_iter17_reg;
            add_i_1_1_3_reg_3327_pp0_iter19_reg <= add_i_1_1_3_reg_3327_pp0_iter18_reg;
            add_i_1_1_3_reg_3327_pp0_iter20_reg <= add_i_1_1_3_reg_3327_pp0_iter19_reg;
            add_i_1_1_3_reg_3327_pp0_iter21_reg <= add_i_1_1_3_reg_3327_pp0_iter20_reg;
            add_i_1_1_3_reg_3327_pp0_iter22_reg <= add_i_1_1_3_reg_3327_pp0_iter21_reg;
            add_i_1_1_3_reg_3327_pp0_iter23_reg <= add_i_1_1_3_reg_3327_pp0_iter22_reg;
            add_i_1_1_3_reg_3327_pp0_iter24_reg <= add_i_1_1_3_reg_3327_pp0_iter23_reg;
            add_i_1_1_3_reg_3327_pp0_iter25_reg <= add_i_1_1_3_reg_3327_pp0_iter24_reg;
            add_i_1_1_3_reg_3327_pp0_iter26_reg <= add_i_1_1_3_reg_3327_pp0_iter25_reg;
            add_i_1_1_3_reg_3327_pp0_iter27_reg <= add_i_1_1_3_reg_3327_pp0_iter26_reg;
            add_i_1_3_3_reg_3391 <= grp_fu_1758_p2;
            add_i_1_3_3_reg_3391_pp0_iter28_reg <= add_i_1_3_3_reg_3391;
            add_i_1_3_3_reg_3391_pp0_iter29_reg <= add_i_1_3_3_reg_3391_pp0_iter28_reg;
            add_i_1_3_3_reg_3391_pp0_iter30_reg <= add_i_1_3_3_reg_3391_pp0_iter29_reg;
            add_i_1_3_3_reg_3391_pp0_iter31_reg <= add_i_1_3_3_reg_3391_pp0_iter30_reg;
            add_i_1_3_3_reg_3391_pp0_iter32_reg <= add_i_1_3_3_reg_3391_pp0_iter31_reg;
            add_i_1_3_3_reg_3391_pp0_iter33_reg <= add_i_1_3_3_reg_3391_pp0_iter32_reg;
            add_i_1_3_3_reg_3391_pp0_iter34_reg <= add_i_1_3_3_reg_3391_pp0_iter33_reg;
            add_i_1_3_3_reg_3391_pp0_iter35_reg <= add_i_1_3_3_reg_3391_pp0_iter34_reg;
            add_i_1_3_3_reg_3391_pp0_iter36_reg <= add_i_1_3_3_reg_3391_pp0_iter35_reg;
            add_i_1_3_3_reg_3391_pp0_iter37_reg <= add_i_1_3_3_reg_3391_pp0_iter36_reg;
            add_i_1_3_3_reg_3391_pp0_iter38_reg <= add_i_1_3_3_reg_3391_pp0_iter37_reg;
            add_i_1_3_3_reg_3391_pp0_iter39_reg <= add_i_1_3_3_reg_3391_pp0_iter38_reg;
            add_i_1_3_3_reg_3391_pp0_iter40_reg <= add_i_1_3_3_reg_3391_pp0_iter39_reg;
            add_i_1_3_3_reg_3391_pp0_iter41_reg <= add_i_1_3_3_reg_3391_pp0_iter40_reg;
            add_i_2_0_3_reg_3333 <= grp_fu_1738_p2;
            add_i_2_0_3_reg_3333_pp0_iter14_reg <= add_i_2_0_3_reg_3333;
            add_i_2_0_3_reg_3333_pp0_iter15_reg <= add_i_2_0_3_reg_3333_pp0_iter14_reg;
            add_i_2_0_3_reg_3333_pp0_iter16_reg <= add_i_2_0_3_reg_3333_pp0_iter15_reg;
            add_i_2_0_3_reg_3333_pp0_iter17_reg <= add_i_2_0_3_reg_3333_pp0_iter16_reg;
            add_i_2_0_3_reg_3333_pp0_iter18_reg <= add_i_2_0_3_reg_3333_pp0_iter17_reg;
            add_i_2_0_3_reg_3333_pp0_iter19_reg <= add_i_2_0_3_reg_3333_pp0_iter18_reg;
            add_i_2_0_3_reg_3333_pp0_iter20_reg <= add_i_2_0_3_reg_3333_pp0_iter19_reg;
            add_i_2_0_3_reg_3333_pp0_iter21_reg <= add_i_2_0_3_reg_3333_pp0_iter20_reg;
            add_i_2_0_3_reg_3333_pp0_iter22_reg <= add_i_2_0_3_reg_3333_pp0_iter21_reg;
            add_i_2_0_3_reg_3333_pp0_iter23_reg <= add_i_2_0_3_reg_3333_pp0_iter22_reg;
            add_i_2_0_3_reg_3333_pp0_iter24_reg <= add_i_2_0_3_reg_3333_pp0_iter23_reg;
            add_i_2_0_3_reg_3333_pp0_iter25_reg <= add_i_2_0_3_reg_3333_pp0_iter24_reg;
            add_i_2_0_3_reg_3333_pp0_iter26_reg <= add_i_2_0_3_reg_3333_pp0_iter25_reg;
            add_i_2_0_3_reg_3333_pp0_iter27_reg <= add_i_2_0_3_reg_3333_pp0_iter26_reg;
            add_i_2_2_3_reg_3340 <= grp_fu_1743_p2;
            add_i_2_2_3_reg_3340_pp0_iter21_reg <= add_i_2_2_3_reg_3340;
            add_i_2_2_3_reg_3340_pp0_iter22_reg <= add_i_2_2_3_reg_3340_pp0_iter21_reg;
            add_i_2_2_3_reg_3340_pp0_iter23_reg <= add_i_2_2_3_reg_3340_pp0_iter22_reg;
            add_i_2_2_3_reg_3340_pp0_iter24_reg <= add_i_2_2_3_reg_3340_pp0_iter23_reg;
            add_i_2_2_3_reg_3340_pp0_iter25_reg <= add_i_2_2_3_reg_3340_pp0_iter24_reg;
            add_i_2_2_3_reg_3340_pp0_iter26_reg <= add_i_2_2_3_reg_3340_pp0_iter25_reg;
            add_i_2_2_3_reg_3340_pp0_iter27_reg <= add_i_2_2_3_reg_3340_pp0_iter26_reg;
            add_i_2_2_3_reg_3340_pp0_iter28_reg <= add_i_2_2_3_reg_3340_pp0_iter27_reg;
            add_i_2_2_3_reg_3340_pp0_iter29_reg <= add_i_2_2_3_reg_3340_pp0_iter28_reg;
            add_i_2_2_3_reg_3340_pp0_iter30_reg <= add_i_2_2_3_reg_3340_pp0_iter29_reg;
            add_i_2_2_3_reg_3340_pp0_iter31_reg <= add_i_2_2_3_reg_3340_pp0_iter30_reg;
            add_i_2_2_3_reg_3340_pp0_iter32_reg <= add_i_2_2_3_reg_3340_pp0_iter31_reg;
            add_i_2_2_3_reg_3340_pp0_iter33_reg <= add_i_2_2_3_reg_3340_pp0_iter32_reg;
            add_i_2_2_3_reg_3340_pp0_iter34_reg <= add_i_2_2_3_reg_3340_pp0_iter33_reg;
            add_i_2_3_3_reg_3397 <= grp_fu_1763_p2;
            add_i_2_3_3_reg_3397_pp0_iter28_reg <= add_i_2_3_3_reg_3397;
            add_i_2_3_3_reg_3397_pp0_iter29_reg <= add_i_2_3_3_reg_3397_pp0_iter28_reg;
            add_i_2_3_3_reg_3397_pp0_iter30_reg <= add_i_2_3_3_reg_3397_pp0_iter29_reg;
            add_i_2_3_3_reg_3397_pp0_iter31_reg <= add_i_2_3_3_reg_3397_pp0_iter30_reg;
            add_i_2_3_3_reg_3397_pp0_iter32_reg <= add_i_2_3_3_reg_3397_pp0_iter31_reg;
            add_i_2_3_3_reg_3397_pp0_iter33_reg <= add_i_2_3_3_reg_3397_pp0_iter32_reg;
            add_i_2_3_3_reg_3397_pp0_iter34_reg <= add_i_2_3_3_reg_3397_pp0_iter33_reg;
            add_i_2_3_3_reg_3397_pp0_iter35_reg <= add_i_2_3_3_reg_3397_pp0_iter34_reg;
            add_i_2_3_3_reg_3397_pp0_iter36_reg <= add_i_2_3_3_reg_3397_pp0_iter35_reg;
            add_i_2_3_3_reg_3397_pp0_iter37_reg <= add_i_2_3_3_reg_3397_pp0_iter36_reg;
            add_i_2_3_3_reg_3397_pp0_iter38_reg <= add_i_2_3_3_reg_3397_pp0_iter37_reg;
            add_i_2_3_3_reg_3397_pp0_iter39_reg <= add_i_2_3_3_reg_3397_pp0_iter38_reg;
            add_i_2_3_3_reg_3397_pp0_iter40_reg <= add_i_2_3_3_reg_3397_pp0_iter39_reg;
            add_i_2_3_3_reg_3397_pp0_iter41_reg <= add_i_2_3_3_reg_3397_pp0_iter40_reg;
            ap_phi_reg_pp0_iter10_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter9_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter10_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter9_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter10_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter9_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter10_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter9_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter10_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter9_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter10_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter9_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter10_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter9_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter10_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter9_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter10_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter9_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter10_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter9_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter10_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter9_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter10_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter9_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter10_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter9_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter10_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter9_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter10_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter9_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter10_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter9_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter10_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter9_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter10_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter9_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter10_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter9_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter10_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter9_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter10_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter9_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter10_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter9_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter10_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter9_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter10_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter9_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter10_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter9_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter10_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter9_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter10_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter9_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter10_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter9_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter10_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter9_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter10_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter9_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter10_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter9_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter10_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter9_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter10_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter9_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter10_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter9_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter10_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter9_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter10_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter9_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter10_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter9_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter10_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter9_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter10_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter9_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter10_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter9_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter10_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter9_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter10_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter9_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter10_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter9_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter10_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter9_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter10_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter9_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter10_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter9_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter10_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter9_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter10_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter9_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter10_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter9_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter10_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter9_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter10_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter9_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter10_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter9_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter10_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter9_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter10_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter9_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter10_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter9_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter10_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter9_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter10_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter9_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter10_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter9_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter10_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter9_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter10_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter9_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter10_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter9_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter10_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter9_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter10_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter9_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter10_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter9_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter11_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter10_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter11_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter10_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter11_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter10_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter11_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter10_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter11_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter10_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter11_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter10_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter11_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter10_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter11_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter10_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter11_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter10_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter11_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter10_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter11_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter10_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter11_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter10_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter11_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter10_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter11_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter10_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter11_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter10_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter11_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter10_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter11_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter10_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter11_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter10_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter11_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter10_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter11_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter10_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter11_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter10_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter11_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter10_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter11_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter10_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter11_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter10_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter11_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter10_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter11_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter10_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter11_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter10_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter11_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter10_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter11_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter10_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter11_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter10_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter11_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter10_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter11_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter10_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter11_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter10_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter11_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter10_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter11_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter10_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter11_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter10_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter11_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter10_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter11_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter10_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter11_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter10_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter11_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter10_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter11_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter10_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter11_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter10_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter11_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter10_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter11_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter10_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter11_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter10_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter11_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter10_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter11_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter10_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter11_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter10_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter11_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter10_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter11_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter10_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter11_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter10_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter11_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter10_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter11_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter10_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter11_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter10_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter11_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter10_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter11_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter10_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter11_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter10_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter11_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter10_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter11_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter10_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter11_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter10_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter11_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter10_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter11_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter10_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter11_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter10_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter11_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter10_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter12_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter11_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter12_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter11_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter12_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter11_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter12_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter11_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter12_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter11_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter12_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter11_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter12_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter11_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter12_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter11_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter12_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter11_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter12_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter11_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter12_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter11_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter12_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter11_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter12_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter11_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter12_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter11_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter12_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter11_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter12_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter11_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter12_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter11_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter12_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter11_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter12_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter11_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter12_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter11_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter12_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter11_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter12_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter11_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter12_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter11_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter12_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter11_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter12_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter11_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter12_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter11_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter12_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter11_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter12_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter11_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter12_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter11_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter12_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter11_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter12_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter11_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter12_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter11_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter12_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter11_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter12_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter11_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter12_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter11_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter12_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter11_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter12_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter11_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter12_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter11_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter12_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter11_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter12_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter11_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter12_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter11_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter12_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter11_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter12_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter11_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter12_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter11_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter12_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter11_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter12_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter11_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter12_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter11_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter12_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter11_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter12_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter11_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter12_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter11_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter12_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter11_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter12_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter11_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter12_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter11_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter12_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter11_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter12_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter11_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter12_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter11_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter12_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter11_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter12_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter11_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter12_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter11_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter12_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter11_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter12_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter11_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter12_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter11_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter12_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter11_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter12_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter11_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter13_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter12_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter13_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter12_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter13_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter12_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter13_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter12_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter13_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter12_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter13_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter12_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter13_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter12_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter13_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter12_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter13_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter12_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter13_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter12_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter13_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter12_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter13_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter12_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter13_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter12_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter13_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter12_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter13_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter12_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter13_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter12_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter13_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter12_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter13_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter12_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter13_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter12_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter13_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter12_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter13_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter12_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter13_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter12_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter13_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter12_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter13_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter12_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter13_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter12_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter13_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter12_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter13_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter12_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter13_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter12_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter13_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter12_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter13_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter12_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter13_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter12_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter13_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter12_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter13_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter12_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter13_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter12_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter13_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter12_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter13_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter12_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter13_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter12_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter13_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter12_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter13_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter12_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter13_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter12_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter13_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter12_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter13_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter12_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter13_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter12_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter13_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter12_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter13_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter12_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter13_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter12_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter13_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter12_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter13_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter12_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter13_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter12_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter13_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter12_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter13_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter12_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter13_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter12_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter13_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter12_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter13_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter12_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter13_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter12_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter13_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter12_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter13_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter12_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter13_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter12_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter13_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter12_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter13_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter12_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter13_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter12_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter13_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter12_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter13_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter12_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter13_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter12_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter14_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter13_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter14_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter13_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter14_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter13_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter14_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter13_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter14_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter13_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter14_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter13_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter14_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter13_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter14_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter13_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter14_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter13_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter14_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter13_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter14_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter13_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter14_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter13_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter14_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter13_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter14_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter13_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter14_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter13_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter14_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter13_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter14_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter13_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter14_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter13_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter14_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter13_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter14_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter13_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter14_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter13_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter14_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter13_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter14_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter13_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter14_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter13_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter14_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter13_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter14_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter13_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter14_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter13_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter14_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter13_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter14_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter13_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter14_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter13_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter14_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter13_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter14_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter13_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter14_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter13_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter14_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter13_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter14_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter13_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter14_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter13_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter14_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter13_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter14_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter13_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter14_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter13_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter14_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter13_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter14_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter13_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter14_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter13_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter14_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter13_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter14_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter13_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter14_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter13_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter14_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter13_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter14_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter13_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter14_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter13_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter14_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter13_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter14_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter13_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter14_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter13_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter14_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter13_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter14_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter13_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter14_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter13_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter14_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter13_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter14_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter13_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter14_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter13_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter14_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter13_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter14_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter13_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter14_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter13_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter14_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter13_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter14_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter13_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter14_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter13_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter14_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter13_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter15_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter14_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter15_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter14_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter15_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter14_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter15_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter14_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter15_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter14_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter15_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter14_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter15_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter14_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter15_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter14_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter15_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter14_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter15_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter14_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter15_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter14_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter15_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter14_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter15_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter14_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter15_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter14_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter15_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter14_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter15_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter14_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter15_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter14_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter15_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter14_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter15_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter14_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter15_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter14_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter15_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter14_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter15_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter14_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter15_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter14_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter15_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter14_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter15_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter14_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter15_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter14_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter15_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter14_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter15_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter14_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter15_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter14_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter15_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter14_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter15_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter14_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter15_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter14_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter15_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter14_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter15_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter14_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter15_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter14_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter15_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter14_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter15_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter14_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter15_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter14_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter15_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter14_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter15_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter14_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter15_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter14_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter15_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter14_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter15_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter14_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter15_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter14_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter15_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter14_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter15_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter14_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter15_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter14_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter15_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter14_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter15_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter14_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter15_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter14_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter15_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter14_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter15_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter14_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter15_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter14_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter15_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter14_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter15_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter14_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter15_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter14_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter15_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter14_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter15_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter14_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter15_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter14_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter15_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter14_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter15_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter14_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter15_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter14_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter15_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter14_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter15_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter14_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter16_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter15_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter16_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter15_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter16_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter15_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter16_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter15_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter16_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter15_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter16_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter15_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter16_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter15_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter16_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter15_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter16_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter15_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter16_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter15_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter16_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter15_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter16_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter15_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter16_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter15_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter16_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter15_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter16_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter15_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter16_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter15_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter16_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter15_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter16_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter15_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter16_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter15_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter16_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter15_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter16_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter15_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter16_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter15_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter16_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter15_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter16_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter15_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter16_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter15_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter16_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter15_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter16_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter15_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter16_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter15_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter16_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter15_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter16_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter15_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter16_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter15_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter16_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter15_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter16_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter15_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter16_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter15_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter16_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter15_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter16_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter15_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter16_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter15_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter16_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter15_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter16_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter15_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter16_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter15_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter16_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter15_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter16_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter15_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter16_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter15_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter16_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter15_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter16_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter15_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter16_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter15_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter16_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter15_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter16_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter15_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter16_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter15_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter16_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter15_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter16_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter15_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter16_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter15_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter16_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter15_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter16_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter15_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter16_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter15_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter16_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter15_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter16_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter15_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter16_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter15_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter16_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter15_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter16_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter15_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter16_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter15_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter16_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter15_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter16_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter15_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter16_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter15_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter17_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter16_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter17_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter16_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter17_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter16_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter17_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter16_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter17_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter16_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter17_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter16_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter17_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter16_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter17_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter16_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter17_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter16_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter17_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter16_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter17_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter16_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter17_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter16_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter17_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter16_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter17_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter16_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter17_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter16_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter17_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter16_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter17_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter16_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter17_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter16_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter17_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter16_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter17_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter16_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter17_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter16_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter17_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter16_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter17_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter16_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter17_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter16_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter17_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter16_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter17_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter16_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter17_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter16_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter17_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter16_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter17_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter16_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter17_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter16_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter17_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter16_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter17_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter16_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter17_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter16_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter17_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter16_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter17_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter16_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter17_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter16_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter17_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter16_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter17_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter16_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter17_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter16_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter17_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter16_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter17_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter16_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter17_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter16_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter17_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter16_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter17_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter16_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter17_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter16_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter17_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter16_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter17_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter16_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter17_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter16_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter17_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter16_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter17_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter16_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter17_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter16_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter17_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter16_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter17_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter16_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter17_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter16_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter17_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter16_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter17_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter16_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter17_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter16_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter17_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter16_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter17_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter16_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter17_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter16_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter17_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter16_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter17_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter16_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter17_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter16_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter17_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter16_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter18_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter17_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter18_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter17_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter18_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter17_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter18_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter17_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter18_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter17_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter18_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter17_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter18_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter17_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter18_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter17_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter18_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter17_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter18_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter17_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter18_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter17_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter18_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter17_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter18_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter17_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter18_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter17_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter18_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter17_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter18_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter17_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter18_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter17_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter18_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter17_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter18_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter17_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter18_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter17_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter18_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter17_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter18_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter17_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter18_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter17_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter18_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter17_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter18_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter17_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter18_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter17_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter18_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter17_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter18_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter17_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter18_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter17_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter18_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter17_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter18_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter17_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter18_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter17_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter18_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter17_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter18_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter17_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter18_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter17_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter18_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter17_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter18_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter17_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter18_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter17_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter18_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter17_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter18_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter17_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter18_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter17_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter18_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter17_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter18_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter17_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter18_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter17_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter18_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter17_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter18_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter17_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter18_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter17_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter18_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter17_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter18_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter17_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter18_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter17_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter18_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter17_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter18_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter17_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter18_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter17_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter18_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter17_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter18_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter17_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter18_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter17_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter18_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter17_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter18_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter17_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter18_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter17_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter18_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter17_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter18_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter17_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter18_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter17_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter18_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter17_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter18_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter17_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter19_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter18_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter19_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter18_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter19_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter18_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter19_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter18_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter19_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter18_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter19_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter18_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter19_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter18_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter19_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter18_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter19_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter18_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter19_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter18_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter19_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter18_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter19_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter18_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter19_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter18_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter19_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter18_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter19_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter18_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter19_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter18_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter19_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter18_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter19_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter18_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter19_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter18_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter19_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter18_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter19_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter18_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter19_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter18_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter19_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter18_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter19_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter18_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter19_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter18_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter19_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter18_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter19_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter18_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter19_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter18_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter19_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter18_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter19_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter18_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter19_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter18_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter19_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter18_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter19_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter18_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter19_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter18_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter19_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter18_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter19_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter18_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter19_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter18_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter19_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter18_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter19_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter18_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter19_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter18_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter19_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter18_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter19_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter18_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter19_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter18_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter19_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter18_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter19_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter18_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter19_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter18_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter19_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter18_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter19_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter18_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter19_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter18_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter19_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter18_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter19_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter18_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter19_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter18_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter19_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter18_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter19_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter18_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter19_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter18_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter19_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter18_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter19_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter18_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter19_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter18_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter19_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter18_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter19_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter18_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter19_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter18_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter19_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter18_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter19_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter18_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter19_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter18_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter20_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter19_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter20_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter19_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter20_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter19_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter20_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter19_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter20_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter19_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter20_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter19_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter20_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter19_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter20_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter19_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter20_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter19_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter20_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter19_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter20_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter19_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter20_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter19_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter20_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter19_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter20_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter19_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter20_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter19_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter20_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter19_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter20_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter19_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter20_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter19_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter20_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter19_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter20_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter19_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter20_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter19_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter20_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter19_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter20_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter19_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter20_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter19_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter20_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter19_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter20_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter19_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter20_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter19_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter20_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter19_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter20_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter19_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter20_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter19_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter20_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter19_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter20_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter19_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter20_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter19_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter20_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter19_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter20_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter19_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter20_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter19_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter20_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter19_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter20_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter19_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter20_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter19_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter20_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter19_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter20_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter19_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter20_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter19_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter20_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter19_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter20_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter19_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter20_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter19_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter20_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter19_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter20_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter19_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter20_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter19_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter20_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter19_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter20_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter19_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter20_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter19_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter20_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter19_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter20_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter19_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter20_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter19_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter20_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter19_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter20_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter19_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter20_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter19_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter20_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter19_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter20_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter19_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter20_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter19_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter20_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter19_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter20_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter19_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter20_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter19_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter20_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter19_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter21_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter20_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter21_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter20_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter21_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter20_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter21_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter20_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter21_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter20_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter21_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter20_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter21_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter20_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter21_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter20_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter21_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter20_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter21_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter20_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter21_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter20_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter21_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter20_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter21_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter20_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter21_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter20_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter21_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter20_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter21_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter20_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter21_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter20_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter21_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter20_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter21_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter20_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter21_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter20_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter21_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter20_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter21_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter20_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter21_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter20_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter21_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter20_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter21_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter20_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter21_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter20_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter21_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter20_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter21_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter20_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter21_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter20_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter21_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter20_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter21_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter20_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter21_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter20_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter21_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter20_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter21_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter20_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter21_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter20_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter21_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter20_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter21_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter20_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter21_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter20_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter21_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter20_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter21_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter20_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter21_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter20_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter21_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter20_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter21_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter20_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter21_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter20_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter21_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter20_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter21_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter20_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter21_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter20_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter21_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter20_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter21_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter20_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter21_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter20_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter21_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter20_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter21_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter20_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter21_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter20_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter21_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter20_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter21_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter20_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter21_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter20_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter21_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter20_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter21_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter20_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter21_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter20_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter21_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter20_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter21_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter20_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter21_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter20_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter21_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter20_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter21_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter20_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter22_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter21_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter22_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter21_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter22_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter21_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter22_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter21_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter22_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter21_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter22_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter21_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter22_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter21_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter22_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter21_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter22_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter21_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter22_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter21_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter22_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter21_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter22_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter21_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter22_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter21_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter22_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter21_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter22_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter21_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter22_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter21_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter22_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter21_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter22_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter21_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter22_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter21_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter22_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter21_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter22_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter21_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter22_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter21_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter22_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter21_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter22_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter21_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter22_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter21_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter22_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter21_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter22_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter21_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter22_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter21_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter22_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter21_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter22_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter21_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter22_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter21_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter22_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter21_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter22_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter21_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter22_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter21_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter22_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter21_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter22_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter21_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter22_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter21_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter22_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter21_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter22_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter21_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter22_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter21_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter22_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter21_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter22_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter21_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter22_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter21_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter22_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter21_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter22_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter21_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter22_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter21_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter22_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter21_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter22_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter21_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter22_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter21_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter22_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter21_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter22_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter21_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter22_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter21_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter22_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter21_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter22_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter21_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter22_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter21_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter22_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter21_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter22_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter21_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter22_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter21_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter22_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter21_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter22_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter21_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter22_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter21_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter22_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter21_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter22_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter21_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter22_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter21_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter23_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter22_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter23_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter22_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter23_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter22_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter23_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter22_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter23_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter22_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter23_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter22_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter23_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter22_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter23_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter22_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter23_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter22_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter23_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter22_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter23_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter22_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter23_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter22_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter23_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter22_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter23_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter22_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter23_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter22_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter23_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter22_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter23_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter22_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter23_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter22_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter23_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter22_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter23_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter22_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter23_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter22_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter23_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter22_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter23_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter22_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter23_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter22_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter23_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter22_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter23_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter22_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter23_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter22_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter23_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter22_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter23_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter22_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter23_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter22_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter23_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter22_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter23_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter22_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter23_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter22_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter23_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter22_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter23_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter22_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter23_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter22_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter23_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter22_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter23_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter22_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter23_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter22_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter23_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter22_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter23_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter22_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter23_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter22_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter23_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter22_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter23_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter22_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter23_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter22_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter23_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter22_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter23_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter22_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter23_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter22_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter23_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter22_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter23_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter22_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter23_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter22_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter23_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter22_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter23_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter22_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter23_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter22_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter23_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter22_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter23_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter22_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter23_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter22_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter23_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter22_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter23_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter22_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter23_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter22_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter23_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter22_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter23_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter22_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter23_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter22_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter23_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter22_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter24_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter23_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter24_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter23_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter24_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter23_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter24_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter23_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter24_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter23_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter24_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter23_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter24_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter23_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter24_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter23_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter24_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter23_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter24_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter23_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter24_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter23_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter24_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter23_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter24_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter23_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter24_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter23_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter24_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter23_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter24_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter23_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter24_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter23_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter24_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter23_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter24_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter23_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter24_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter23_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter24_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter23_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter24_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter23_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter24_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter23_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter24_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter23_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter24_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter23_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter24_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter23_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter24_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter23_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter24_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter23_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter24_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter23_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter24_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter23_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter24_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter23_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter24_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter23_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter24_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter23_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter24_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter23_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter24_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter23_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter24_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter23_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter24_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter23_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter24_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter23_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter24_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter23_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter24_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter23_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter24_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter23_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter24_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter23_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter24_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter23_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter24_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter23_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter24_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter23_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter24_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter23_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter24_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter23_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter24_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter23_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter24_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter23_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter24_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter23_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter24_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter23_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter24_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter23_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter24_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter23_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter24_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter23_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter24_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter23_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter24_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter23_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter24_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter23_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter24_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter23_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter24_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter23_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter24_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter23_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter24_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter23_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter24_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter23_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter24_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter23_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter24_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter23_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter25_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter24_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter25_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter24_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter25_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter24_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter25_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter24_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter25_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter24_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter25_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter24_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter25_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter24_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter25_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter24_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter25_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter24_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter25_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter24_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter25_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter24_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter25_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter24_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter25_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter24_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter25_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter24_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter25_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter24_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter25_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter24_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter25_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter24_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter25_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter24_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter25_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter24_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter25_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter24_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter25_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter24_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter25_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter24_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter25_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter24_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter25_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter24_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter25_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter24_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter25_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter24_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter25_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter24_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter25_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter24_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter25_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter24_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter25_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter24_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter25_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter24_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter25_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter24_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter25_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter24_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter25_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter24_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter25_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter24_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter25_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter24_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter25_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter24_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter25_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter24_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter25_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter24_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter25_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter24_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter25_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter24_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter25_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter24_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter25_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter24_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter25_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter24_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter25_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter24_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter25_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter24_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter25_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter24_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter25_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter24_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter25_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter24_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter25_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter24_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter25_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter24_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter25_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter24_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter25_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter24_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter25_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter24_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter25_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter24_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter25_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter24_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter25_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter24_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter25_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter24_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter25_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter24_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter25_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter24_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter25_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter24_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter25_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter24_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter25_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter24_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter25_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter24_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter26_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter25_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter26_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter25_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter26_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter25_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter26_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter25_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter26_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter25_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter26_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter25_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter26_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter25_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter26_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter25_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter26_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter25_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter26_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter25_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter26_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter25_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter26_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter25_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter26_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter25_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter26_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter25_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter26_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter25_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter26_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter25_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter26_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter25_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter26_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter25_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter26_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter25_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter26_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter25_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter26_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter25_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter26_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter25_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter26_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter25_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter26_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter25_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter26_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter25_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter26_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter25_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter26_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter25_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter26_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter25_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter26_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter25_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter26_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter25_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter26_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter25_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter26_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter25_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter26_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter25_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter26_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter25_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter26_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter25_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter26_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter25_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter26_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter25_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter26_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter25_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter26_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter25_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter26_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter25_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter26_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter25_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter26_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter25_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter26_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter25_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter26_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter25_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter26_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter25_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter26_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter25_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter26_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter25_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter26_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter25_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter26_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter25_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter26_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter25_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter26_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter25_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter26_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter25_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter26_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter25_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter26_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter25_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter26_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter25_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter26_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter25_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter26_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter25_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter26_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter25_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter26_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter25_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter26_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter25_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter26_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter25_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter26_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter25_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter26_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter25_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter26_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter25_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter27_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter26_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter27_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter26_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter27_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter26_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter27_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter26_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter27_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter26_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter27_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter26_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter27_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter26_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter27_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter26_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter27_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter26_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter27_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter26_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter27_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter26_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter27_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter26_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter27_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter26_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter27_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter26_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter27_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter26_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter27_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter26_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter27_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter26_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter27_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter26_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter27_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter26_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter27_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter26_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter27_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter26_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter27_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter26_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter27_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter26_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter27_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter26_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter27_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter26_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter27_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter26_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter27_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter26_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter27_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter26_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter27_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter26_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter27_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter26_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter27_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter26_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter27_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter26_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter27_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter26_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter27_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter26_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter27_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter26_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter27_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter26_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter27_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter26_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter27_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter26_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter27_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter26_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter27_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter26_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter27_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter26_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter27_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter26_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter27_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter26_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter27_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter26_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter27_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter26_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter27_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter26_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter27_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter26_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter27_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter26_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter27_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter26_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter27_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter26_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter27_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter26_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter27_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter26_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter27_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter26_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter27_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter26_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter27_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter26_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter27_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter26_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter27_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter26_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter27_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter26_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter27_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter26_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter27_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter26_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter27_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter26_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter27_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter26_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter27_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter26_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter27_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter26_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter28_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter27_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter28_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter27_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter28_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter27_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter28_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter27_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter28_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter27_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter28_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter27_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter28_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter27_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter28_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter27_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter28_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter27_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter28_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter27_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter28_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter27_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter28_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter27_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter28_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter27_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter28_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter27_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter28_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter27_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter28_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter27_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter28_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter27_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter28_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter27_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter28_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter27_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter28_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter27_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter28_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter27_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter28_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter27_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter28_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter27_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter28_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter27_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter28_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter27_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter28_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter27_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter28_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter27_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter28_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter27_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter28_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter27_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter28_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter27_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter28_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter27_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter28_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter27_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter28_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter27_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter28_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter27_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter28_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter27_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter28_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter27_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter28_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter27_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter28_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter27_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter28_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter27_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter28_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter27_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter28_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter27_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter28_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter27_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter28_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter27_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter28_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter27_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter28_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter27_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter28_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter27_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter28_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter27_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter28_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter27_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter28_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter27_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter28_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter27_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter28_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter27_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter28_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter27_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter28_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter27_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter28_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter27_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter28_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter27_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter28_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter27_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter28_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter27_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter28_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter27_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter28_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter27_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter28_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter27_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter28_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter27_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter28_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter27_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter28_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter27_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter28_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter27_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter29_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter28_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter29_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter28_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter29_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter28_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter29_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter28_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter29_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter28_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter29_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter28_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter29_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter28_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter29_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter28_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter29_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter28_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter29_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter28_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter29_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter28_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter29_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter28_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter29_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter28_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter29_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter28_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter29_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter28_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter29_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter28_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter29_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter28_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter29_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter28_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter29_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter28_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter29_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter28_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter29_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter28_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter29_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter28_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter29_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter28_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter29_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter28_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter29_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter28_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter29_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter28_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter29_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter28_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter29_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter28_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter29_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter28_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter29_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter28_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter29_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter28_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter29_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter28_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter29_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter28_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter29_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter28_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter29_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter28_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter29_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter28_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter29_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter28_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter29_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter28_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter29_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter28_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter29_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter28_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter29_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter28_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter29_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter28_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter29_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter28_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter29_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter28_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter29_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter28_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter29_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter28_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter29_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter28_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter29_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter28_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter29_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter28_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter29_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter28_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter29_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter28_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter29_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter28_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter29_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter28_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter29_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter28_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter29_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter28_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter29_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter28_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter29_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter28_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter29_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter28_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter29_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter28_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter29_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter28_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter29_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter28_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter29_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter28_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter29_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter28_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter29_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter28_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter2_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter1_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter2_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter1_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter2_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter1_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter2_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter1_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter2_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter1_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter2_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter1_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter2_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter1_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter2_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter1_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter2_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter1_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter2_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter1_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter2_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter1_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter2_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter1_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter2_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter1_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter2_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter1_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter2_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter1_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter2_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter1_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter2_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter1_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter2_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter1_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter2_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter1_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter2_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter1_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter2_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter1_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter2_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter1_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter2_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter1_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter2_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter1_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter2_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter1_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter2_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter1_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter2_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter1_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter2_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter1_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter2_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter1_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter2_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter1_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter2_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter1_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter2_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter1_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter2_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter1_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter2_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter1_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter2_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter1_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter2_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter1_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter2_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter1_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter2_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter1_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter2_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter1_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter2_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter1_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter2_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter1_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter2_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter1_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter2_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter1_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter2_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter1_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter2_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter1_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter2_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter1_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter2_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter1_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter2_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter1_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter2_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter1_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter2_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter1_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter2_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter1_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter2_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter1_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter2_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter1_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter2_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter1_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter2_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter1_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter2_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter1_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter2_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter1_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter2_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter1_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter2_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter1_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter2_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter1_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter2_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter1_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter2_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter1_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter2_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter1_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter2_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter1_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter30_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter29_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter30_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter29_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter30_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter29_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter30_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter29_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter30_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter29_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter30_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter29_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter30_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter29_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter30_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter29_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter30_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter29_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter30_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter29_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter30_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter29_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter30_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter29_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter30_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter29_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter30_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter29_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter30_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter29_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter30_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter29_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter30_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter29_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter30_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter29_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter30_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter29_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter30_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter29_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter30_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter29_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter30_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter29_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter30_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter29_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter30_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter29_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter30_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter29_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter30_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter29_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter30_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter29_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter30_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter29_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter30_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter29_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter30_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter29_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter30_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter29_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter30_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter29_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter30_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter29_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter30_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter29_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter30_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter29_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter30_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter29_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter30_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter29_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter30_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter29_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter30_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter29_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter30_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter29_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter30_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter29_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter30_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter29_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter30_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter29_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter30_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter29_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter30_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter29_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter30_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter29_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter30_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter29_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter30_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter29_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter30_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter29_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter30_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter29_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter30_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter29_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter30_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter29_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter30_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter29_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter30_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter29_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter30_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter29_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter30_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter29_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter30_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter29_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter30_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter29_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter30_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter29_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter30_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter29_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter30_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter29_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter30_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter29_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter30_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter29_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter30_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter29_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter31_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter30_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter31_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter30_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter31_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter30_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter31_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter30_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter31_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter30_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter31_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter30_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter31_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter30_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter31_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter30_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter31_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter30_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter31_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter30_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter31_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter30_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter31_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter30_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter31_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter30_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter31_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter30_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter31_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter30_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter31_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter30_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter31_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter30_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter31_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter30_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter31_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter30_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter31_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter30_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter31_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter30_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter31_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter30_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter31_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter30_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter31_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter30_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter31_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter30_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter31_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter30_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter31_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter30_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter31_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter30_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter31_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter30_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter31_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter30_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter31_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter30_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter31_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter30_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter31_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter30_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter31_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter30_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter31_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter30_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter31_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter30_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter31_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter30_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter31_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter30_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter31_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter30_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter31_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter30_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter31_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter30_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter31_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter30_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter31_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter30_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter31_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter30_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter31_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter30_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter31_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter30_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter31_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter30_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter31_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter30_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter31_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter30_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter31_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter30_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter31_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter30_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter31_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter30_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter31_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter30_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter31_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter30_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter31_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter30_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter31_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter30_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter31_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter30_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter31_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter30_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter31_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter30_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter31_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter30_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter31_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter30_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter31_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter30_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter31_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter30_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter31_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter30_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter32_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter31_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter32_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter31_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter32_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter31_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter32_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter31_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter32_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter31_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter32_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter31_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter32_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter31_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter32_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter31_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter32_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter31_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter32_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter31_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter32_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter31_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter32_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter31_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter32_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter31_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter32_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter31_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter32_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter31_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter32_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter31_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter32_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter31_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter32_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter31_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter32_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter31_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter32_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter31_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter32_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter31_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter32_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter31_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter32_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter31_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter32_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter31_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter32_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter31_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter32_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter31_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter32_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter31_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter32_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter31_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter32_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter31_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter32_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter31_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter32_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter31_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter32_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter31_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter32_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter31_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter32_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter31_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter32_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter31_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter32_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter31_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter32_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter31_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter32_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter31_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter32_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter31_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter32_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter31_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter32_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter31_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter32_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter31_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter32_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter31_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter32_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter31_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter32_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter31_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter32_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter31_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter32_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter31_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter32_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter31_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter32_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter31_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter32_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter31_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter32_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter31_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter32_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter31_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter32_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter31_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter32_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter31_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter32_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter31_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter32_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter31_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter32_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter31_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter32_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter31_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter32_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter31_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter32_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter31_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter32_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter31_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter32_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter31_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter32_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter31_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter32_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter31_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter33_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter32_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter33_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter32_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter33_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter32_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter33_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter32_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter33_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter32_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter33_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter32_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter33_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter32_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter33_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter32_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter33_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter32_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter33_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter32_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter33_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter32_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter33_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter32_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter33_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter32_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter33_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter32_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter33_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter32_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter33_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter32_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter33_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter32_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter33_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter32_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter33_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter32_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter33_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter32_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter33_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter32_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter33_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter32_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter33_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter32_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter33_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter32_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter33_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter32_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter33_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter32_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter33_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter32_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter33_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter32_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter33_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter32_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter33_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter32_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter33_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter32_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter33_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter32_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter33_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter32_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter33_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter32_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter33_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter32_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter33_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter32_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter33_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter32_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter33_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter32_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter33_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter32_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter33_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter32_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter33_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter32_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter33_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter32_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter33_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter32_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter33_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter32_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter33_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter32_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter33_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter32_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter33_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter32_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter33_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter32_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter33_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter32_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter33_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter32_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter33_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter32_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter33_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter32_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter33_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter32_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter33_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter32_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter33_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter32_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter33_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter32_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter33_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter32_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter33_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter32_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter33_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter32_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter33_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter32_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter33_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter32_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter33_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter32_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter33_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter32_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter33_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter32_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter34_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter33_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter34_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter33_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter34_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter33_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter34_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter33_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter34_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter33_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter34_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter33_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter34_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter33_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter34_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter33_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter34_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter33_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter34_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter33_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter34_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter33_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter34_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter33_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter34_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter33_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter34_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter33_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter34_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter33_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter34_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter33_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter34_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter33_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter34_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter33_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter34_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter33_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter34_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter33_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter34_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter33_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter34_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter33_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter34_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter33_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter34_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter33_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter34_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter33_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter34_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter33_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter34_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter33_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter34_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter33_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter34_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter33_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter34_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter33_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter34_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter33_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter34_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter33_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter34_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter33_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter34_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter33_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter34_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter33_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter34_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter33_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter34_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter33_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter34_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter33_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter34_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter33_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter34_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter33_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter34_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter33_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter34_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter33_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter34_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter33_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter34_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter33_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter34_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter33_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter34_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter33_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter34_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter33_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter34_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter33_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter34_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter33_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter34_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter33_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter34_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter33_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter34_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter33_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter34_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter33_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter34_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter33_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter34_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter33_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter34_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter33_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter34_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter33_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter34_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter33_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter34_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter33_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter34_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter33_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter34_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter33_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter34_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter33_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter34_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter33_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter34_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter33_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter35_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter34_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter35_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter34_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter35_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter34_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter35_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter34_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter35_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter34_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter35_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter34_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter35_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter34_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter35_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter34_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter35_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter34_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter35_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter34_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter35_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter34_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter35_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter34_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter35_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter34_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter35_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter34_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter35_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter34_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter35_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter34_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter35_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter34_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter35_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter34_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter35_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter34_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter35_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter34_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter35_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter34_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter35_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter34_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter35_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter34_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter35_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter34_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter35_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter34_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter35_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter34_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter35_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter34_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter35_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter34_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter35_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter34_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter35_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter34_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter35_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter34_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter35_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter34_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter35_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter34_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter35_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter34_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter35_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter34_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter35_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter34_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter35_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter34_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter35_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter34_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter35_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter34_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter35_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter34_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter35_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter34_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter35_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter34_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter35_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter34_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter35_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter34_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter35_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter34_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter35_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter34_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter35_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter34_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter35_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter34_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter35_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter34_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter35_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter34_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter35_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter34_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter35_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter34_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter35_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter34_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter35_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter34_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter35_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter34_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter35_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter34_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter35_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter34_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter35_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter34_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter35_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter34_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter35_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter34_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter35_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter34_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter35_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter34_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter35_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter34_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter35_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter34_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter36_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter35_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter36_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter35_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter36_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter35_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter36_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter35_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter36_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter35_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter36_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter35_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter36_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter35_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter36_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter35_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter36_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter35_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter36_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter35_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter36_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter35_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter36_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter35_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter36_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter35_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter36_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter35_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter36_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter35_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter36_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter35_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter36_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter35_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter36_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter35_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter36_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter35_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter36_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter35_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter36_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter35_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter36_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter35_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter36_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter35_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter36_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter35_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter36_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter35_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter36_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter35_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter36_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter35_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter36_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter35_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter36_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter35_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter36_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter35_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter36_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter35_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter36_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter35_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter36_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter35_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter36_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter35_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter36_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter35_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter36_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter35_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter36_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter35_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter36_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter35_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter36_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter35_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter36_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter35_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter36_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter35_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter36_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter35_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter36_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter35_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter36_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter35_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter36_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter35_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter36_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter35_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter36_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter35_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter36_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter35_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter36_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter35_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter36_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter35_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter36_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter35_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter36_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter35_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter36_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter35_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter36_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter35_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter36_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter35_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter36_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter35_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter36_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter35_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter36_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter35_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter36_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter35_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter36_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter35_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter36_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter35_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter36_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter35_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter36_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter35_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter36_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter35_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter37_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter36_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter37_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter36_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter37_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter36_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter37_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter36_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter37_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter36_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter37_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter36_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter37_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter36_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter37_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter36_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter37_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter36_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter37_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter36_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter37_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter36_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter37_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter36_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter37_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter36_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter37_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter36_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter37_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter36_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter37_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter36_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter37_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter36_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter37_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter36_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter37_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter36_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter37_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter36_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter37_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter36_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter37_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter36_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter37_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter36_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter37_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter36_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter37_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter36_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter37_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter36_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter37_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter36_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter37_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter36_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter37_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter36_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter37_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter36_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter37_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter36_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter37_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter36_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter37_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter36_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter37_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter36_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter37_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter36_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter37_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter36_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter37_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter36_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter37_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter36_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter37_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter36_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter37_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter36_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter37_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter36_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter37_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter36_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter37_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter36_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter37_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter36_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter37_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter36_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter37_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter36_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter37_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter36_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter37_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter36_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter37_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter36_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter37_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter36_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter37_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter36_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter37_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter36_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter37_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter36_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter37_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter36_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter37_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter36_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter37_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter36_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter37_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter36_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter37_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter36_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter37_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter36_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter37_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter36_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter37_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter36_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter37_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter36_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter37_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter36_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter37_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter36_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter38_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter37_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter38_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter37_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter38_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter37_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter38_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter37_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter38_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter37_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter38_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter37_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter38_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter37_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter38_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter37_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter38_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter37_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter38_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter37_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter38_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter37_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter38_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter37_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter38_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter37_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter38_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter37_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter38_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter37_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter38_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter37_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter38_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter37_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter38_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter37_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter38_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter37_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter38_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter37_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter38_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter37_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter38_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter37_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter38_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter37_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter38_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter37_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter38_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter37_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter38_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter37_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter38_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter37_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter38_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter37_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter38_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter37_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter38_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter37_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter38_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter37_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter38_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter37_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter38_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter37_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter38_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter37_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter38_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter37_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter38_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter37_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter38_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter37_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter38_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter37_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter38_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter37_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter38_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter37_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter38_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter37_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter38_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter37_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter38_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter37_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter38_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter37_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter38_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter37_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter38_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter37_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter38_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter37_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter38_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter37_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter38_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter37_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter38_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter37_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter38_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter37_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter38_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter37_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter38_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter37_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter38_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter37_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter38_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter37_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter38_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter37_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter38_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter37_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter38_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter37_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter38_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter37_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter38_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter37_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter38_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter37_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter38_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter37_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter38_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter37_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter38_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter37_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter39_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter38_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter39_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter38_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter39_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter38_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter39_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter38_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter39_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter38_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter39_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter38_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter39_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter38_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter39_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter38_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter39_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter38_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter39_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter38_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter39_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter38_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter39_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter38_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter39_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter38_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter39_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter38_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter39_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter38_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter39_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter38_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter39_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter38_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter39_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter38_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter39_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter38_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter39_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter38_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter39_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter38_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter39_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter38_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter39_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter38_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter39_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter38_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter39_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter38_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter39_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter38_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter39_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter38_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter39_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter38_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter39_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter38_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter39_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter38_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter39_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter38_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter39_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter38_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter39_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter38_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter39_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter38_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter39_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter38_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter39_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter38_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter39_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter38_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter39_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter38_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter39_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter38_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter39_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter38_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter39_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter38_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter39_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter38_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter39_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter38_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter39_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter38_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter39_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter38_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter39_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter38_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter39_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter38_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter39_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter38_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter39_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter38_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter39_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter38_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter39_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter38_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter39_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter38_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter39_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter38_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter39_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter38_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter39_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter38_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter39_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter38_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter39_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter38_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter39_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter38_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter39_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter38_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter39_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter38_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter39_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter38_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter39_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter38_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter39_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter38_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter39_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter38_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter3_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter2_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter3_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter2_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter3_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter2_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter3_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter2_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter3_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter2_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter3_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter2_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter3_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter2_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter3_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter2_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter3_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter2_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter3_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter2_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter3_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter2_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter3_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter2_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter3_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter2_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter3_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter2_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter3_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter2_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter3_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter2_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter3_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter2_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter3_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter2_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter3_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter2_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter3_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter2_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter3_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter2_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter3_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter2_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter3_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter2_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter3_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter2_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter3_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter2_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter3_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter2_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter3_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter2_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter3_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter2_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter3_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter2_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter3_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter2_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter3_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter2_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter3_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter2_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter3_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter2_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter3_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter2_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter3_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter2_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter3_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter2_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter3_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter2_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter3_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter2_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter3_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter2_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter3_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter2_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter3_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter2_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter3_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter2_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter3_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter2_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter3_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter2_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter3_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter2_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter3_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter2_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter3_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter2_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter3_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter2_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter3_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter2_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter3_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter2_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter3_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter2_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter3_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter2_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter3_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter2_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter3_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter2_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter3_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter2_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter3_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter2_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter3_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter2_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter3_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter2_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter3_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter2_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter3_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter2_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter3_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter2_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter3_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter2_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter3_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter2_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter3_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter2_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter40_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter39_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter40_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter39_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter40_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter39_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter40_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter39_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter40_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter39_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter40_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter39_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter40_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter39_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter40_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter39_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter40_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter39_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter40_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter39_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter40_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter39_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter40_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter39_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter40_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter39_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter40_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter39_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter40_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter39_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter40_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter39_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter40_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter39_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter40_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter39_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter40_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter39_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter40_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter39_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter40_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter39_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter40_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter39_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter40_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter39_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter40_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter39_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter40_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter39_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter40_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter39_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter40_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter39_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter40_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter39_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter40_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter39_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter40_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter39_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter40_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter39_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter40_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter39_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter40_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter39_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter40_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter39_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter40_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter39_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter40_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter39_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter40_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter39_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter40_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter39_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter40_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter39_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter40_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter39_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter40_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter39_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter40_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter39_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter40_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter39_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter40_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter39_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter40_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter39_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter40_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter39_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter40_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter39_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter40_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter39_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter40_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter39_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter40_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter39_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter40_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter39_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter40_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter39_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter40_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter39_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter40_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter39_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter40_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter39_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter40_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter39_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter40_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter39_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter40_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter39_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter40_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter39_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter40_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter39_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter40_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter39_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter40_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter39_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter40_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter39_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter40_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter39_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter41_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter40_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter41_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter40_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter41_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter40_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter41_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter40_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter41_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter40_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter41_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter40_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter41_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter40_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter41_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter40_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter41_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter40_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter41_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter40_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter41_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter40_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter41_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter40_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter41_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter40_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter41_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter40_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter41_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter40_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter41_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter40_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter41_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter40_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter41_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter40_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter41_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter40_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter41_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter40_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter41_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter40_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter41_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter40_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter41_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter40_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter41_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter40_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter41_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter40_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter41_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter40_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter41_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter40_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter41_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter40_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter41_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter40_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter41_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter40_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter41_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter40_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter41_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter40_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter41_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter40_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter41_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter40_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter41_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter40_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter41_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter40_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter41_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter40_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter41_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter40_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter41_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter40_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter41_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter40_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter41_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter40_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter41_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter40_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter41_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter40_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter41_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter40_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter41_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter40_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter41_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter40_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter41_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter40_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter41_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter40_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter41_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter40_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter41_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter40_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter41_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter40_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter41_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter40_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter41_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter40_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter41_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter40_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter41_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter40_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter41_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter40_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter41_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter40_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter41_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter40_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter41_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter40_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter41_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter40_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter41_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter40_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter41_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter40_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter41_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter40_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter41_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter40_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter42_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter41_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter42_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter41_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter42_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter41_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter42_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter41_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter42_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter41_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter42_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter41_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter42_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter41_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter42_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter41_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter42_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter41_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter42_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter41_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter42_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter41_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter42_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter41_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter42_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter41_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter42_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter41_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter42_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter41_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter42_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter41_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter42_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter41_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter42_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter41_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter42_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter41_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter42_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter41_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter42_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter41_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter42_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter41_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter42_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter41_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter42_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter41_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter42_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter41_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter42_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter41_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter42_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter41_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter42_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter41_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter42_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter41_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter42_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter41_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter42_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter41_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter42_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter41_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter42_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter41_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter42_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter41_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter42_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter41_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter42_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter41_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter42_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter41_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter42_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter41_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter42_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter41_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter42_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter41_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter42_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter41_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter42_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter41_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter42_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter41_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter42_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter41_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter42_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter41_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter42_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter41_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter42_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter41_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter42_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter41_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter42_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter41_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter42_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter41_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter42_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter41_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter42_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter41_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter42_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter41_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter42_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter41_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter42_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter41_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter42_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter41_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter42_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter41_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter42_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter41_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter42_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter41_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter42_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter41_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter42_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter41_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter42_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter41_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter42_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter41_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter42_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter41_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter43_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter42_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter43_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter42_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter43_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter42_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter43_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter42_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter43_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter42_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter43_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter42_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter43_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter42_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter43_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter42_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter43_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter42_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter43_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter42_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter43_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter42_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter43_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter42_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter43_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter42_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter43_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter42_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter43_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter42_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter43_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter42_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter43_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter42_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter43_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter42_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter43_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter42_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter43_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter42_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter43_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter42_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter43_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter42_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter43_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter42_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter43_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter42_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter43_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter42_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter43_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter42_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter43_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter42_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter43_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter42_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter43_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter42_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter43_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter42_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter43_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter42_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter43_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter42_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter43_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter42_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter43_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter42_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter43_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter42_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter43_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter42_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter43_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter42_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter43_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter42_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter43_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter42_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter43_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter42_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter43_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter42_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter43_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter42_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter43_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter42_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter43_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter42_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter43_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter42_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter43_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter42_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter43_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter42_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter43_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter42_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter43_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter42_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter43_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter42_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter43_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter42_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter43_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter42_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter43_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter42_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter43_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter42_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter43_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter42_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter43_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter42_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter43_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter42_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter43_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter42_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter43_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter42_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter43_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter42_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter43_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter42_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter43_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter42_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter43_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter42_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter43_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter42_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter44_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter43_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter44_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter43_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter44_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter43_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter44_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter43_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter44_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter43_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter44_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter43_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter44_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter43_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter44_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter43_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter44_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter43_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter44_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter43_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter44_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter43_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter44_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter43_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter44_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter43_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter44_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter43_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter44_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter43_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter44_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter43_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter44_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter43_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter44_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter43_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter44_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter43_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter44_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter43_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter44_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter43_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter44_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter43_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter44_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter43_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter44_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter43_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter44_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter43_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter44_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter43_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter44_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter43_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter44_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter43_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter44_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter43_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter44_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter43_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter44_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter43_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter44_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter43_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter44_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter43_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter44_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter43_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter44_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter43_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter44_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter43_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter44_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter43_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter44_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter43_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter44_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter43_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter44_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter43_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter44_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter43_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter44_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter43_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter44_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter43_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter44_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter43_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter44_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter43_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter44_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter43_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter44_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter43_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter44_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter43_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter44_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter43_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter44_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter43_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter44_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter43_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter44_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter43_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter44_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter43_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter44_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter43_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter44_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter43_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter44_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter43_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter44_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter43_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter44_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter43_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter44_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter43_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter44_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter43_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter44_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter43_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter44_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter43_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter44_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter43_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter44_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter43_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter45_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter44_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter45_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter44_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter45_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter44_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter45_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter44_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter45_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter44_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter45_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter44_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter45_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter44_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter45_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter44_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter45_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter44_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter45_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter44_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter45_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter44_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter45_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter44_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter45_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter44_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter45_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter44_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter45_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter44_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter45_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter44_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter45_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter44_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter45_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter44_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter45_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter44_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter45_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter44_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter45_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter44_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter45_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter44_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter45_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter44_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter45_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter44_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter45_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter44_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter45_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter44_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter45_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter44_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter45_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter44_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter45_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter44_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter45_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter44_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter45_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter44_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter45_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter44_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter45_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter44_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter45_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter44_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter45_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter44_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter45_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter44_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter45_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter44_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter45_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter44_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter45_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter44_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter45_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter44_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter45_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter44_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter45_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter44_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter45_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter44_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter45_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter44_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter45_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter44_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter45_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter44_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter45_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter44_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter45_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter44_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter45_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter44_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter45_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter44_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter45_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter44_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter45_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter44_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter45_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter44_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter45_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter44_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter45_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter44_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter45_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter44_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter45_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter44_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter45_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter44_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter45_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter44_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter45_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter44_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter45_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter44_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter45_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter44_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter45_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter44_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter45_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter44_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter46_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter45_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter46_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter45_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter46_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter45_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter46_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter45_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter46_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter45_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter46_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter45_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter46_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter45_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter46_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter45_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter46_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter45_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter46_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter45_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter46_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter45_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter46_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter45_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter46_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter45_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter46_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter45_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter46_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter45_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter46_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter45_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter46_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter45_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter46_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter45_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter46_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter45_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter46_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter45_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter46_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter45_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter46_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter45_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter46_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter45_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter46_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter45_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter46_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter45_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter46_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter45_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter46_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter45_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter46_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter45_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter46_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter45_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter46_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter45_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter46_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter45_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter46_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter45_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter46_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter45_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter46_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter45_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter46_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter45_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter46_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter45_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter46_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter45_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter46_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter45_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter46_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter45_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter46_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter45_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter46_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter45_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter46_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter45_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter46_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter45_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter46_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter45_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter46_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter45_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter46_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter45_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter46_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter45_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter46_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter45_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter46_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter45_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter46_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter45_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter46_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter45_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter46_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter45_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter46_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter45_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter46_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter45_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter46_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter45_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter46_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter45_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter46_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter45_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter46_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter45_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter46_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter45_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter46_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter45_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter46_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter45_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter46_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter45_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter46_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter45_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter46_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter45_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter47_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter46_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter47_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter46_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter47_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter46_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter47_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter46_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter47_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter46_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter47_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter46_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter47_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter46_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter47_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter46_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter47_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter46_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter47_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter46_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter47_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter46_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter47_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter46_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter47_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter46_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter47_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter46_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter47_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter46_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter47_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter46_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter47_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter46_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter47_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter46_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter47_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter46_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter47_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter46_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter47_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter46_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter47_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter46_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter47_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter46_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter47_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter46_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter47_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter46_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter47_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter46_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter47_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter46_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter47_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter46_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter47_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter46_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter47_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter46_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter47_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter46_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter47_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter46_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter47_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter46_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter47_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter46_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter47_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter46_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter47_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter46_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter47_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter46_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter47_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter46_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter47_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter46_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter47_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter46_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter47_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter46_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter47_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter46_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter47_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter46_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter47_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter46_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter47_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter46_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter47_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter46_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter47_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter46_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter47_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter46_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter47_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter46_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter47_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter46_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter47_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter46_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter47_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter46_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter47_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter46_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter47_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter46_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter47_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter46_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter47_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter46_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter47_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter46_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter47_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter46_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter47_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter46_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter47_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter46_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter47_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter46_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter47_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter46_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter47_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter46_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter47_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter46_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter48_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter47_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter48_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter47_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter48_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter47_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter48_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter47_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter48_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter47_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter48_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter47_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter48_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter47_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter48_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter47_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter48_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter47_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter48_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter47_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter48_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter47_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter48_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter47_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter48_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter47_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter48_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter47_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter48_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter47_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter48_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter47_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter48_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter47_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter48_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter47_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter48_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter47_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter48_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter47_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter48_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter47_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter48_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter47_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter48_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter47_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter48_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter47_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter48_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter47_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter48_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter47_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter48_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter47_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter48_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter47_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter48_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter47_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter48_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter47_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter48_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter47_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter48_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter47_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter48_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter47_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter48_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter47_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter48_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter47_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter48_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter47_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter48_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter47_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter48_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter47_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter48_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter47_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter48_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter47_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter48_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter47_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter48_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter47_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter48_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter47_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter48_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter47_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter48_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter47_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter48_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter47_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter48_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter47_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter48_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter47_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter48_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter47_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter48_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter47_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter48_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter47_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter48_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter47_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter48_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter47_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter48_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter47_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter48_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter47_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter48_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter47_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter48_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter47_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter48_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter47_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter48_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter47_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter48_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter47_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter48_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter47_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter48_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter47_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter48_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter47_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter48_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter47_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter49_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter48_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter49_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter48_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter49_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter48_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter49_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter48_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter49_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter48_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter49_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter48_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter49_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter48_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter49_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter48_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter49_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter48_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter49_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter48_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter49_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter48_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter49_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter48_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter49_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter48_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter49_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter48_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter49_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter48_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter49_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter48_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter49_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter48_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter49_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter48_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter49_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter48_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter49_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter48_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter49_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter48_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter49_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter48_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter49_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter48_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter49_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter48_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter49_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter48_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter49_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter48_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter49_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter48_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter49_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter48_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter49_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter48_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter49_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter48_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter49_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter48_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter49_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter48_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter49_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter48_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter49_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter48_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter49_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter48_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter49_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter48_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter49_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter48_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter49_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter48_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter49_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter48_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter49_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter48_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter49_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter48_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter49_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter48_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter49_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter48_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter49_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter48_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter49_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter48_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter49_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter48_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter49_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter48_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter49_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter48_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter49_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter48_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter49_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter48_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter49_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter48_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter49_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter48_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter49_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter48_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter49_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter48_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter49_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter48_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter49_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter48_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter49_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter48_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter49_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter48_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter49_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter48_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter49_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter48_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter49_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter48_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter49_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter48_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter49_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter48_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter49_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter48_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter4_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter3_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter4_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter3_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter4_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter3_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter4_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter3_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter4_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter3_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter4_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter3_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter4_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter3_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter4_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter3_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter4_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter3_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter4_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter3_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter4_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter3_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter4_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter3_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter4_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter3_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter4_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter3_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter4_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter3_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter4_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter3_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter4_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter3_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter4_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter3_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter4_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter3_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter4_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter3_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter4_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter3_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter4_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter3_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter4_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter3_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter4_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter3_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter4_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter3_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter4_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter3_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter4_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter3_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter4_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter3_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter4_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter3_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter4_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter3_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter4_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter3_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter4_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter3_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter4_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter3_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter4_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter3_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter4_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter3_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter4_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter3_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter4_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter3_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter4_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter3_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter4_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter3_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter4_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter3_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter4_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter3_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter4_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter3_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter4_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter3_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter4_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter3_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter4_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter3_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter4_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter3_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter4_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter3_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter4_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter3_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter4_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter3_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter4_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter3_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter4_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter3_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter4_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter3_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter4_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter3_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter4_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter3_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter4_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter3_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter4_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter3_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter4_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter3_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter4_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter3_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter4_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter3_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter4_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter3_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter4_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter3_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter4_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter3_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter4_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter3_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter4_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter3_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter50_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter49_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter50_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter49_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter50_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter49_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter50_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter49_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter50_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter49_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter50_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter49_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter50_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter49_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter50_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter49_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter50_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter49_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter50_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter49_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter50_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter49_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter50_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter49_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter50_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter49_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter50_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter49_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter50_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter49_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter50_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter49_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter50_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter49_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter50_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter49_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter50_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter49_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter50_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter49_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter50_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter49_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter50_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter49_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter50_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter49_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter50_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter49_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter50_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter49_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter50_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter49_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter50_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter49_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter50_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter49_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter50_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter49_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter50_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter49_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter50_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter49_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter50_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter49_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter50_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter49_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter50_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter49_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter50_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter49_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter50_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter49_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter50_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter49_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter50_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter49_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter50_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter49_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter50_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter49_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter50_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter49_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter50_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter49_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter50_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter49_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter50_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter49_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter50_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter49_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter50_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter49_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter50_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter49_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter50_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter49_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter50_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter49_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter50_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter49_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter50_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter49_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter50_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter49_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter50_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter49_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter50_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter49_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter50_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter49_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter50_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter49_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter50_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter49_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter50_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter49_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter50_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter49_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter50_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter49_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter50_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter49_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter50_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter49_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter50_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter49_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter50_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter49_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter51_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter50_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter51_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter50_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter51_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter50_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter51_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter50_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter51_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter50_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter51_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter50_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter51_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter50_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter51_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter50_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter51_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter50_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter51_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter50_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter51_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter50_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter51_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter50_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter51_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter50_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter51_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter50_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter51_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter50_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter51_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter50_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter51_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter50_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter51_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter50_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter51_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter50_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter51_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter50_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter51_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter50_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter51_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter50_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter51_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter50_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter51_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter50_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter51_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter50_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter51_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter50_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter51_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter50_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter51_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter50_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter51_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter50_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter51_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter50_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter51_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter50_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter51_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter50_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter51_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter50_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter51_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter50_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter51_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter50_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter51_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter50_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter51_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter50_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter51_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter50_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter51_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter50_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter51_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter50_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter51_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter50_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter51_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter50_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter51_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter50_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter51_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter50_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter51_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter50_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter51_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter50_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter51_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter50_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter51_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter50_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter51_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter50_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter51_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter50_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter51_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter50_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter51_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter50_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter51_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter50_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter51_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter50_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter51_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter50_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter51_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter50_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter51_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter50_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter51_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter50_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter51_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter50_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter51_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter50_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter51_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter50_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter51_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter50_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter51_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter50_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter51_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter50_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter52_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter51_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter52_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter51_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter52_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter51_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter52_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter51_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter52_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter51_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter52_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter51_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter52_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter51_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter52_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter51_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter52_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter51_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter52_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter51_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter52_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter51_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter52_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter51_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter52_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter51_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter52_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter51_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter52_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter51_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter52_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter51_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter52_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter51_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter52_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter51_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter52_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter51_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter52_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter51_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter52_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter51_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter52_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter51_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter52_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter51_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter52_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter51_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter52_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter51_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter52_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter51_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter52_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter51_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter52_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter51_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter52_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter51_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter52_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter51_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter52_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter51_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter52_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter51_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter52_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter51_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter52_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter51_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter52_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter51_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter52_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter51_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter52_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter51_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter52_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter51_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter52_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter51_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter52_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter51_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter52_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter51_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter52_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter51_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter52_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter51_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter52_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter51_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter52_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter51_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter52_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter51_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter52_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter51_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter52_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter51_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter52_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter51_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter52_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter51_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter52_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter51_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter52_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter51_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter52_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter51_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter52_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter51_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter52_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter51_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter52_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter51_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter52_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter51_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter52_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter51_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter52_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter51_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter52_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter51_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter52_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter51_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter52_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter51_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter52_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter51_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter52_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter51_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter53_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter52_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter53_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter52_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter53_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter52_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter53_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter52_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter53_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter52_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter53_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter52_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter53_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter52_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter53_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter52_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter53_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter52_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter53_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter52_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter53_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter52_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter53_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter52_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter53_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter52_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter53_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter52_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter53_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter52_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter53_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter52_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter53_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter52_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter53_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter52_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter53_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter52_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter53_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter52_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter53_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter52_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter53_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter52_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter53_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter52_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter53_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter52_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter53_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter52_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter53_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter52_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter53_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter52_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter53_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter52_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter53_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter52_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter53_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter52_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter53_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter52_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter53_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter52_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter53_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter52_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter53_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter52_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter53_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter52_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter53_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter52_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter53_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter52_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter53_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter52_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter53_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter52_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter53_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter52_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter53_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter52_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter53_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter52_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter53_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter52_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter53_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter52_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter53_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter52_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter53_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter52_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter53_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter52_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter53_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter52_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter53_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter52_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter53_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter52_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter53_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter52_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter53_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter52_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter53_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter52_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter53_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter52_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter53_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter52_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter53_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter52_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter53_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter52_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter53_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter52_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter53_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter52_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter53_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter52_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter53_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter52_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter53_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter52_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter53_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter52_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter53_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter52_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter54_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter53_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter54_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter53_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter54_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter53_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter54_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter53_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter54_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter53_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter54_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter53_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter54_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter53_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter54_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter53_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter54_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter53_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter54_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter53_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter54_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter53_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter54_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter53_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter54_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter53_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter54_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter53_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter54_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter53_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter54_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter53_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter54_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter53_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter54_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter53_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter54_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter53_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter54_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter53_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter54_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter53_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter54_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter53_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter54_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter53_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter54_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter53_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter54_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter53_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter54_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter53_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter54_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter53_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter54_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter53_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter54_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter53_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter54_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter53_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter54_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter53_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter54_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter53_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter54_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter53_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter54_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter53_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter54_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter53_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter54_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter53_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter54_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter53_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter54_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter53_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter54_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter53_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter54_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter53_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter54_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter53_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter54_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter53_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter54_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter53_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter54_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter53_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter54_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter53_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter54_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter53_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter54_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter53_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter54_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter53_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter54_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter53_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter54_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter53_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter54_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter53_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter54_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter53_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter54_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter53_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter54_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter53_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter54_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter53_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter54_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter53_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter54_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter53_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter54_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter53_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter54_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter53_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter54_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter53_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter54_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter53_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter54_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter53_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter54_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter53_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter54_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter53_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter55_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter54_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter55_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter54_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter55_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter54_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter55_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter54_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter55_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter54_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter55_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter54_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter55_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter54_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter55_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter54_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter55_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter54_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter55_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter54_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter55_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter54_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter55_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter54_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter55_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter54_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter55_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter54_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter55_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter54_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter55_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter54_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter55_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter54_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter55_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter54_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter55_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter54_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter55_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter54_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter55_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter54_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter55_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter54_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter55_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter54_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter55_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter54_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter55_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter54_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter55_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter54_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter55_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter54_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter55_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter54_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter55_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter54_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter55_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter54_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter55_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter54_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter55_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter54_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter55_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter54_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter55_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter54_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter55_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter54_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter55_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter54_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter55_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter54_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter55_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter54_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter55_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter54_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter55_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter54_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter55_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter54_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter55_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter54_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter55_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter54_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter55_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter54_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter55_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter54_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter55_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter54_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter55_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter54_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter55_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter54_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter55_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter54_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter55_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter54_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter55_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter54_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter55_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter54_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter55_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter54_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter55_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter54_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter55_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter54_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter55_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter54_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter55_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter54_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter55_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter54_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter55_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter54_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter55_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter54_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter55_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter54_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter55_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter54_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter55_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter54_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter55_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter54_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter56_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter55_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter56_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter55_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter56_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter55_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter56_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter55_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter56_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter55_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter56_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter55_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter56_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter55_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter56_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter55_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter56_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter55_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter56_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter55_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter56_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter55_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter56_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter55_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter56_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter55_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter56_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter55_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter56_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter55_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter56_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter55_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter56_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter55_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter56_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter55_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter56_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter55_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter56_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter55_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter56_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter55_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter56_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter55_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter56_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter55_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter56_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter55_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter56_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter55_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter56_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter55_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter56_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter55_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter56_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter55_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter56_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter55_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter56_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter55_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter56_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter55_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter56_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter55_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter56_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter55_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter56_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter55_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter56_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter55_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter56_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter55_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter56_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter55_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter56_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter55_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter56_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter55_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter56_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter55_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter56_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter55_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter56_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter55_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter56_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter55_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter56_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter55_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter56_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter55_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter56_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter55_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter56_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter55_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter56_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter55_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter56_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter55_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter56_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter55_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter56_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter55_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter56_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter55_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter56_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter55_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter56_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter55_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter56_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter55_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter56_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter55_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter56_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter55_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter56_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter55_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter56_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter55_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter56_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter55_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter56_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter55_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter56_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter55_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter56_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter55_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter56_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter55_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter57_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter56_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter57_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter56_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter57_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter56_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter57_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter56_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter57_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter56_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter57_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter56_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter57_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter56_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter57_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter56_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter57_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter56_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter57_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter56_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter57_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter56_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter57_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter56_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter57_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter56_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter57_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter56_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter57_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter56_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter57_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter56_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter57_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter56_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter57_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter56_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter57_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter56_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter57_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter56_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter57_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter56_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter57_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter56_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter57_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter56_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter57_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter56_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter57_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter56_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter57_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter56_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter57_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter56_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter57_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter56_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter57_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter56_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter57_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter56_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter57_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter56_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter57_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter56_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter57_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter56_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter57_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter56_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter57_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter56_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter57_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter56_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter57_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter56_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter57_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter56_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter57_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter56_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter57_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter56_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter57_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter56_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter57_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter56_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter57_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter56_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter57_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter56_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter57_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter56_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter57_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter56_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter57_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter56_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter57_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter56_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter57_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter56_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter57_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter56_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter57_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter56_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter57_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter56_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter57_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter56_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter57_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter56_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter57_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter56_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter57_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter56_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter57_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter56_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter57_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter56_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter57_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter56_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter57_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter56_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter57_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter56_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter57_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter56_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter57_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter56_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter57_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter56_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter58_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter57_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter58_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter57_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter58_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter57_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter58_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter57_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter58_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter57_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter58_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter57_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter58_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter57_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter58_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter57_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter58_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter57_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter58_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter57_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter58_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter57_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter58_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter57_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter58_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter57_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter58_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter57_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter58_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter57_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter58_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter57_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter58_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter57_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter58_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter57_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter58_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter57_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter58_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter57_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter58_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter57_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter58_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter57_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter58_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter57_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter58_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter57_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter58_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter57_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter58_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter57_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter58_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter57_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter58_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter57_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter58_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter57_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter58_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter57_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter58_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter57_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter58_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter57_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter58_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter57_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter58_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter57_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter58_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter57_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter58_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter57_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter58_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter57_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter58_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter57_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter58_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter57_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter58_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter57_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter58_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter57_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter58_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter57_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter58_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter57_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter58_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter57_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter58_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter57_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter58_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter57_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter58_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter57_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter58_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter57_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter58_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter57_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter58_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter57_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter58_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter57_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter58_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter57_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter58_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter57_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter58_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter57_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter58_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter57_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter58_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter57_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter58_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter57_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter58_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter57_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter58_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter57_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter58_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter57_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter58_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter57_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter58_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter57_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter58_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter57_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter58_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter57_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter59_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter58_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter59_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter58_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter59_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter58_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter59_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter58_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter59_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter58_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter59_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter58_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter59_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter58_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter59_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter58_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter59_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter58_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter59_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter58_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter59_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter58_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter59_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter58_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter59_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter58_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter59_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter58_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter59_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter58_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter59_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter58_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter59_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter58_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter59_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter58_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter59_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter58_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter59_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter58_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter59_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter58_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter59_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter58_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter59_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter58_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter59_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter58_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter59_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter58_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter59_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter58_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter59_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter58_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter59_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter58_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter59_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter58_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter59_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter58_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter59_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter58_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter59_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter58_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter59_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter58_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter59_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter58_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter59_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter58_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter59_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter58_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter59_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter58_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter59_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter58_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter59_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter58_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter59_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter58_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter59_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter58_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter59_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter58_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter59_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter58_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter59_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter58_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter59_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter58_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter59_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter58_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter59_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter58_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter59_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter58_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter59_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter58_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter59_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter58_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter59_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter58_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter59_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter58_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter59_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter58_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter59_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter58_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter59_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter58_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter59_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter58_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter59_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter58_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter59_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter58_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter59_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter58_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter59_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter58_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter59_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter58_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter59_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter58_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter59_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter58_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter59_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter58_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter5_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter4_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter5_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter4_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter5_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter4_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter5_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter4_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter5_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter4_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter5_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter4_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter5_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter4_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter5_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter4_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter5_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter4_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter5_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter4_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter5_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter4_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter5_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter4_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter5_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter4_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter5_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter4_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter5_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter4_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter5_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter4_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter5_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter4_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter5_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter4_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter5_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter4_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter5_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter4_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter5_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter4_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter5_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter4_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter5_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter4_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter5_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter4_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter5_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter4_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter5_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter4_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter5_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter4_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter5_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter4_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter5_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter4_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter5_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter4_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter5_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter4_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter5_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter4_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter5_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter4_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter5_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter4_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter5_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter4_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter5_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter4_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter5_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter4_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter5_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter4_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter5_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter4_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter5_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter4_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter5_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter4_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter5_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter4_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter5_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter4_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter5_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter4_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter5_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter4_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter5_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter4_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter5_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter4_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter5_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter4_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter5_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter4_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter5_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter4_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter5_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter4_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter5_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter4_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter5_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter4_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter5_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter4_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter5_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter4_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter5_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter4_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter5_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter4_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter5_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter4_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter5_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter4_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter5_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter4_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter5_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter4_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter5_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter4_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter5_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter4_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter5_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter4_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter60_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter59_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter60_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter59_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter60_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter59_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter60_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter59_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter60_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter59_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter60_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter59_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter60_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter59_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter60_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter59_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter60_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter59_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter60_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter59_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter60_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter59_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter60_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter59_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter60_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter59_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter60_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter59_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter60_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter59_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter60_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter59_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter60_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter59_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter60_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter59_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter60_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter59_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter60_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter59_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter60_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter59_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter60_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter59_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter60_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter59_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter60_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter59_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter60_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter59_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter60_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter59_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter60_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter59_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter60_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter59_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter60_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter59_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter60_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter59_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter60_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter59_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter60_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter59_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter60_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter59_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter60_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter59_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter60_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter59_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter60_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter59_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter60_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter59_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter60_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter59_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter60_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter59_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter60_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter59_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter60_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter59_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter60_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter59_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter60_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter59_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter60_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter59_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter60_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter59_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter60_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter59_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter60_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter59_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter60_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter59_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter60_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter59_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter60_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter59_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter60_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter59_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter60_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter59_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter60_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter59_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter60_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter59_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter60_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter59_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter60_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter59_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter60_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter59_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter60_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter59_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter60_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter59_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter60_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter59_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter60_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter59_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter60_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter59_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter60_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter59_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter60_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter59_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter61_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter60_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter61_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter60_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter61_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter60_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter61_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter60_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter61_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter60_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter61_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter60_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter61_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter60_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter61_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter60_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter61_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter60_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter61_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter60_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter61_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter60_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter61_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter60_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter61_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter60_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter61_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter60_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter61_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter60_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter61_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter60_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter61_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter60_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter61_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter60_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter61_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter60_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter61_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter60_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter61_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter60_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter61_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter60_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter61_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter60_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter61_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter60_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter61_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter60_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter61_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter60_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter61_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter60_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter61_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter60_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter61_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter60_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter61_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter60_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter61_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter60_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter61_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter60_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter61_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter60_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter61_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter60_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter61_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter60_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter61_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter60_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter61_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter60_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter61_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter60_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter61_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter60_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter61_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter60_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter61_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter60_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter61_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter60_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter61_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter60_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter61_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter60_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter61_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter60_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter61_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter60_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter61_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter60_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter61_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter60_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter61_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter60_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter61_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter60_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter61_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter60_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter61_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter60_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter61_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter60_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter61_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter60_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter61_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter60_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter61_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter60_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter61_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter60_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter61_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter60_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter61_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter60_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter61_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter60_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter61_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter60_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter61_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter60_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter61_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter60_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter61_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter60_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter62_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter61_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter62_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter61_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter62_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter61_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter62_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter61_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter62_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter61_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter62_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter61_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter62_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter61_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter62_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter61_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter62_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter61_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter62_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter61_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter62_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter61_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter62_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter61_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter62_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter61_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter62_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter61_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter62_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter61_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter62_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter61_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter62_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter61_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter62_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter61_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter62_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter61_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter62_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter61_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter62_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter61_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter62_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter61_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter62_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter61_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter62_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter61_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter62_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter61_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter62_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter61_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter62_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter61_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter62_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter61_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter62_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter61_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter62_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter61_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter62_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter61_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter62_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter61_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter62_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter61_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter62_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter61_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter62_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter61_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter62_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter61_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter62_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter61_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter62_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter61_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter62_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter61_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter62_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter61_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter62_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter61_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter62_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter61_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter62_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter61_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter62_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter61_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter62_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter61_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter62_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter61_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter62_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter61_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter62_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter61_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter62_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter61_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter62_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter61_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter62_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter61_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter62_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter61_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter62_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter61_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter62_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter61_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter62_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter61_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter62_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter61_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter62_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter61_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter62_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter61_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter62_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter61_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter62_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter61_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter62_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter61_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter62_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter61_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter62_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter61_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter62_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter61_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter63_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter62_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter63_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter62_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter63_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter62_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter63_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter62_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter63_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter62_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter63_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter62_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter63_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter62_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter63_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter62_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter63_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter62_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter63_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter62_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter63_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter62_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter63_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter62_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter63_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter62_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter63_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter62_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter63_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter62_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter63_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter62_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter63_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter62_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter63_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter62_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter63_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter62_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter63_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter62_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter63_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter62_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter63_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter62_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter63_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter62_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter63_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter62_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter63_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter62_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter63_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter62_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter63_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter62_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter63_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter62_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter63_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter62_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter63_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter62_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter63_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter62_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter63_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter62_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter63_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter62_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter63_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter62_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter63_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter62_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter63_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter62_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter63_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter62_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter63_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter62_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter63_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter62_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter63_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter62_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter63_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter62_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter63_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter62_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter63_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter62_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter63_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter62_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter63_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter62_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter63_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter62_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter63_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter62_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter63_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter62_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter63_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter62_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter63_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter62_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter63_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter62_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter63_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter62_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter63_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter62_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter63_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter62_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter63_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter62_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter63_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter62_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter63_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter62_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter63_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter62_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter63_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter62_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter63_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter62_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter63_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter62_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter63_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter62_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter63_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter62_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter63_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter62_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter64_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter63_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter64_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter63_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter64_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter63_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter64_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter63_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter64_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter63_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter64_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter63_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter64_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter63_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter64_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter63_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter64_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter63_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter64_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter63_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter64_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter63_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter64_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter63_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter64_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter63_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter64_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter63_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter64_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter63_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter64_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter63_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter64_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter63_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter64_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter63_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter64_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter63_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter64_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter63_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter64_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter63_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter64_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter63_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter64_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter63_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter64_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter63_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter64_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter63_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter64_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter63_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter64_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter63_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter64_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter63_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter64_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter63_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter64_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter63_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter64_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter63_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter64_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter63_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter64_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter63_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter64_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter63_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter64_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter63_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter64_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter63_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter64_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter63_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter64_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter63_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter64_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter63_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter64_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter63_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter64_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter63_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter64_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter63_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter64_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter63_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter64_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter63_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter64_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter63_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter64_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter63_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter64_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter63_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter64_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter63_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter64_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter63_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter64_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter63_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter64_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter63_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter64_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter63_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter64_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter63_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter64_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter63_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter64_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter63_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter64_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter63_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter64_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter63_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter64_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter63_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter64_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter63_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter64_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter63_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter64_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter63_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter64_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter63_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter64_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter63_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter64_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter63_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter65_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter64_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter65_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter64_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter65_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter64_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter65_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter64_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter65_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter64_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter65_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter64_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter65_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter64_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter65_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter64_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter65_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter64_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter65_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter64_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter65_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter64_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter65_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter64_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter65_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter64_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter65_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter64_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter65_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter64_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter65_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter64_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter65_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter64_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter65_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter64_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter65_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter64_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter65_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter64_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter65_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter64_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter65_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter64_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter65_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter64_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter65_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter64_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter65_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter64_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter65_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter64_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter65_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter64_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter65_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter64_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter65_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter64_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter65_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter64_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter65_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter64_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter65_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter64_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter65_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter64_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter65_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter64_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter65_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter64_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter65_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter64_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter65_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter64_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter65_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter64_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter65_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter64_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter65_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter64_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter65_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter64_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter65_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter64_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter65_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter64_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter65_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter64_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter65_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter64_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter65_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter64_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter65_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter64_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter65_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter64_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter65_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter64_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter65_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter64_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter65_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter64_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter65_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter64_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter65_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter64_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter65_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter64_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter65_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter64_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter65_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter64_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter65_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter64_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter65_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter64_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter65_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter64_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter65_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter64_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter65_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter64_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter65_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter64_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter65_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter64_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter65_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter64_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter66_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter65_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter66_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter65_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter66_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter65_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter66_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter65_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter66_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter65_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter66_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter65_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter66_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter65_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter66_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter65_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter66_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter65_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter66_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter65_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter66_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter65_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter66_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter65_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter66_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter65_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter66_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter65_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter66_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter65_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter66_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter65_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter66_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter65_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter66_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter65_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter66_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter65_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter66_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter65_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter66_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter65_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter66_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter65_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter66_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter65_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter66_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter65_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter66_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter65_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter66_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter65_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter66_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter65_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter66_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter65_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter66_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter65_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter66_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter65_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter66_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter65_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter66_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter65_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter66_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter65_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter66_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter65_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter66_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter65_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter66_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter65_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter66_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter65_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter66_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter65_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter66_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter65_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter66_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter65_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter66_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter65_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter66_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter65_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter66_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter65_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter66_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter65_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter66_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter65_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter66_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter65_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter66_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter65_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter66_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter65_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter66_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter65_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter66_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter65_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter66_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter65_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter66_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter65_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter66_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter65_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter66_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter65_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter66_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter65_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter66_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter65_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter66_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter65_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter66_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter65_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter66_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter65_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter66_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter65_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter66_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter65_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter66_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter65_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter66_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter65_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter66_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter65_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter67_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter66_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter67_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter66_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter67_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter66_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter67_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter66_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter67_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter66_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter67_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter66_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter67_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter66_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter67_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter66_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter67_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter66_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter67_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter66_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter67_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter66_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter67_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter66_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter67_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter66_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter67_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter66_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter67_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter66_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter67_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter66_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter67_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter66_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter67_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter66_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter67_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter66_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter67_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter66_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter67_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter66_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter67_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter66_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter67_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter66_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter67_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter66_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter67_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter66_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter67_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter66_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter67_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter66_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter67_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter66_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter67_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter66_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter67_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter66_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter67_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter66_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter67_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter66_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter67_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter66_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter67_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter66_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter67_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter66_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter67_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter66_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter67_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter66_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter67_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter66_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter67_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter66_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter67_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter66_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter67_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter66_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter67_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter66_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter67_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter66_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter67_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter66_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter67_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter66_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter67_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter66_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter67_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter66_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter67_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter66_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter67_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter66_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter67_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter66_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter67_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter66_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter67_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter66_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter67_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter66_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter67_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter66_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter67_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter66_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter67_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter66_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter67_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter66_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter67_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter66_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter67_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter66_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter67_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter66_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter67_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter66_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter67_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter66_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter67_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter66_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter67_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter66_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter68_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter67_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter68_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter67_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter68_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter67_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter68_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter67_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter68_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter67_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter68_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter67_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter68_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter67_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter68_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter67_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter68_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter67_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter68_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter67_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter68_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter67_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter68_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter67_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter68_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter67_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter68_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter67_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter68_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter67_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter68_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter67_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter68_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter67_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter68_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter67_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter68_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter67_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter68_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter67_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter68_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter67_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter68_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter67_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter68_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter67_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter68_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter67_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter68_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter67_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter68_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter67_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter68_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter67_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter68_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter67_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter68_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter67_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter68_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter67_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter68_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter67_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter68_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter67_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter68_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter67_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter68_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter67_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter68_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter67_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter68_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter67_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter68_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter67_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter68_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter67_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter68_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter67_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter68_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter67_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter68_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter67_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter68_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter67_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter68_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter67_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter68_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter67_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter68_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter67_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter68_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter67_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter68_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter67_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter68_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter67_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter68_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter67_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter68_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter67_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter68_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter67_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter68_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter67_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter68_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter67_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter68_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter67_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter68_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter67_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter68_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter67_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter68_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter67_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter68_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter67_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter68_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter67_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter68_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter67_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter68_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter67_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter68_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter67_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter68_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter67_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter68_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter67_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter69_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter68_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter69_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter68_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter69_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter68_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter69_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter68_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter69_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter68_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter69_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter68_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter69_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter68_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter69_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter68_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter69_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter68_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter69_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter68_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter69_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter68_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter69_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter68_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter69_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter68_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter69_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter68_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter69_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter68_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter69_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter68_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter69_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter68_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter69_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter68_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter69_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter68_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter69_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter68_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter69_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter68_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter69_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter68_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter69_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter68_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter69_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter68_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter69_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter68_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter69_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter68_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter69_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter68_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter69_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter68_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter69_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter68_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter69_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter68_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter69_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter68_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter69_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter68_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter69_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter68_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter69_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter68_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter69_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter68_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter69_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter68_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter69_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter68_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter69_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter68_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter69_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter68_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter69_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter68_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter69_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter68_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter69_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter68_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter69_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter68_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter69_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter68_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter69_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter68_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter69_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter68_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter69_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter68_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter69_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter68_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter69_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter68_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter69_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter68_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter69_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter68_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter69_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter68_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter69_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter68_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter69_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter68_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter69_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter68_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter69_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter68_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter69_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter68_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter69_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter68_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter69_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter68_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter69_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter68_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter69_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter68_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter69_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter68_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter69_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter68_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter69_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter68_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter6_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter5_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter6_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter5_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter6_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter5_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter6_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter5_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter6_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter5_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter6_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter5_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter6_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter5_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter6_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter5_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter6_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter5_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter6_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter5_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter6_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter5_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter6_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter5_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter6_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter5_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter6_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter5_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter6_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter5_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter6_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter5_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter6_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter5_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter6_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter5_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter6_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter5_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter6_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter5_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter6_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter5_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter6_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter5_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter6_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter5_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter6_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter5_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter6_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter5_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter6_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter5_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter6_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter5_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter6_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter5_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter6_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter5_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter6_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter5_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter6_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter5_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter6_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter5_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter6_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter5_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter6_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter5_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter6_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter5_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter6_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter5_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter6_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter5_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter6_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter5_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter6_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter5_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter6_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter5_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter6_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter5_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter6_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter5_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter6_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter5_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter6_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter5_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter6_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter5_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter6_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter5_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter6_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter5_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter6_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter5_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter6_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter5_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter6_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter5_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter6_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter5_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter6_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter5_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter6_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter5_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter6_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter5_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter6_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter5_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter6_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter5_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter6_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter5_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter6_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter5_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter6_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter5_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter6_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter5_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter6_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter5_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter6_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter5_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter6_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter5_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter6_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter5_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter70_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter69_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter70_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter69_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter70_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter69_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter70_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter69_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter70_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter69_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter70_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter69_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter70_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter69_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter70_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter69_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter70_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter69_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter70_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter69_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter70_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter69_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter70_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter69_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter70_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter69_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter70_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter69_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter70_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter69_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter70_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter69_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter70_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter69_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter70_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter69_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter70_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter69_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter70_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter69_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter70_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter69_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter70_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter69_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter70_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter69_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter70_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter69_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter70_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter69_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter70_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter69_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter70_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter69_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter70_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter69_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter70_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter69_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter70_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter69_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter70_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter69_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter70_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter69_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter70_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter69_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter70_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter69_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter70_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter69_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter70_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter69_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter70_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter69_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter70_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter69_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter70_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter69_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter70_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter69_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter70_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter69_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter70_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter69_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter70_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter69_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter70_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter69_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter70_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter69_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter70_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter69_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter70_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter69_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter70_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter69_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter70_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter69_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter70_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter69_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter70_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter69_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter70_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter69_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter70_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter69_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter70_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter69_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter70_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter69_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter70_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter69_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter70_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter69_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter70_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter69_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter70_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter69_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter70_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter69_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter70_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter69_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter70_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter69_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter70_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter69_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter70_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter69_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter71_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter70_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter71_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter70_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter71_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter70_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter71_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter70_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter71_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter70_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter71_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter70_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter71_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter70_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter71_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter70_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter71_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter70_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter71_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter70_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter71_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter70_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter71_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter70_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter71_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter70_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter71_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter70_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter71_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter70_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter71_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter70_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter71_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter70_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter71_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter70_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter71_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter70_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter71_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter70_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter71_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter70_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter71_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter70_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter71_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter70_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter71_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter70_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter71_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter70_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter71_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter70_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter71_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter70_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter71_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter70_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter71_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter70_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter71_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter70_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter71_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter70_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter71_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter70_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter71_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter70_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter71_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter70_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter71_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter70_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter71_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter70_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter71_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter70_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter71_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter70_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter71_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter70_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter71_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter70_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter71_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter70_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter71_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter70_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter71_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter70_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter71_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter70_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter71_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter70_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter71_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter70_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter71_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter70_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter71_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter70_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter71_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter70_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter71_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter70_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter71_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter70_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter71_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter70_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter71_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter70_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter71_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter70_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter71_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter70_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter71_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter70_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter71_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter70_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter71_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter70_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter71_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter70_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter71_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter70_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter71_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter70_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter71_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter70_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter71_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter70_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter71_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter70_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter72_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter71_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter72_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter71_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter72_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter71_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter72_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter71_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter72_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter71_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter72_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter71_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter72_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter71_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter72_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter71_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter72_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter71_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter72_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter71_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter72_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter71_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter72_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter71_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter72_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter71_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter72_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter71_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter72_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter71_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter72_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter71_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter72_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter71_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter72_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter71_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter72_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter71_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter72_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter71_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter72_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter71_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter72_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter71_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter72_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter71_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter72_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter71_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter72_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter71_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter72_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter71_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter72_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter71_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter72_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter71_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter72_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter71_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter72_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter71_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter72_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter71_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter72_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter71_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter72_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter71_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter72_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter71_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter72_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter71_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter72_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter71_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter72_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter71_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter72_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter71_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter72_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter71_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter72_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter71_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter72_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter71_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter72_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter71_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter72_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter71_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter72_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter71_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter72_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter71_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter72_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter71_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter72_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter71_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter72_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter71_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter72_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter71_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter72_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter71_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter72_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter71_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter72_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter71_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter72_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter71_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter72_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter71_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter72_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter71_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter72_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter71_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter72_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter71_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter72_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter71_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter72_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter71_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter72_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter71_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter72_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter71_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter72_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter71_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter72_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter71_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter72_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter71_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter73_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter72_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter73_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter72_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter73_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter72_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter73_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter72_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter73_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter72_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter73_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter72_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter73_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter72_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter73_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter72_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter73_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter72_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter73_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter72_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter73_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter72_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter73_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter72_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter73_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter72_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter73_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter72_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter73_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter72_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter73_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter72_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter73_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter72_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter73_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter72_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter73_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter72_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter73_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter72_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter73_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter72_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter73_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter72_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter73_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter72_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter73_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter72_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter73_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter72_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter73_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter72_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter73_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter72_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter73_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter72_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter73_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter72_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter73_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter72_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter73_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter72_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter73_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter72_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter73_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter72_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter73_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter72_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter73_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter72_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter73_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter72_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter73_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter72_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter73_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter72_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter73_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter72_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter73_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter72_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter73_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter72_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter73_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter72_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter73_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter72_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter73_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter72_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter73_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter72_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter73_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter72_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter73_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter72_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter73_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter72_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter73_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter72_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter73_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter72_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter73_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter72_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter73_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter72_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter73_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter72_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter73_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter72_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter73_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter72_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter73_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter72_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter73_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter72_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter73_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter72_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter73_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter72_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter73_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter72_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter73_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter72_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter73_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter72_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter73_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter72_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter73_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter72_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter74_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter73_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter74_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter73_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter74_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter73_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter74_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter73_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter74_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter73_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter74_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter73_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter74_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter73_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter74_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter73_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter74_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter73_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter74_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter73_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter74_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter73_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter74_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter73_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter74_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter73_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter74_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter73_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter74_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter73_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter74_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter73_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter74_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter73_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter74_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter73_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter74_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter73_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter74_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter73_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter74_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter73_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter74_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter73_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter74_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter73_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter74_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter73_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter74_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter73_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter74_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter73_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter74_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter73_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter74_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter73_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter74_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter73_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter74_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter73_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter74_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter73_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter74_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter73_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter74_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter73_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter74_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter73_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter74_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter73_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter74_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter73_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter74_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter73_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter74_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter73_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter74_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter73_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter74_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter73_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter74_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter73_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter74_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter73_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter74_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter73_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter74_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter73_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter74_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter73_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter74_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter73_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter74_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter73_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter74_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter73_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter74_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter73_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter74_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter73_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter74_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter73_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter74_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter73_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter74_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter73_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter74_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter73_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter74_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter73_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter74_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter73_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter74_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter73_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter74_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter73_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter74_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter73_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter74_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter73_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter74_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter73_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter74_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter73_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter74_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter73_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter74_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter73_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter75_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter74_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter75_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter74_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter75_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter74_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter75_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter74_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter75_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter74_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter75_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter74_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter75_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter74_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter75_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter74_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter75_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter74_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter75_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter74_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter75_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter74_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter75_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter74_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter75_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter74_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter75_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter74_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter75_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter74_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter75_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter74_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter75_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter74_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter75_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter74_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter75_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter74_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter75_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter74_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter75_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter74_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter75_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter74_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter75_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter74_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter75_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter74_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter75_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter74_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter75_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter74_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter75_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter74_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter75_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter74_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter75_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter74_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter75_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter74_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter75_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter74_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter75_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter74_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter75_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter74_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter75_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter74_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter75_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter74_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter75_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter74_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter75_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter74_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter75_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter74_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter75_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter74_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter75_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter74_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter75_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter74_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter75_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter74_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter75_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter74_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter75_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter74_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter75_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter74_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter75_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter74_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter75_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter74_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter75_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter74_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter75_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter74_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter75_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter74_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter75_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter74_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter75_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter74_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter75_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter74_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter75_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter74_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter75_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter74_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter75_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter74_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter75_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter74_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter75_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter74_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter75_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter74_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter75_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter74_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter75_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter74_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter75_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter74_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter75_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter74_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter75_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter74_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter76_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter75_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter76_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter75_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter76_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter75_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter76_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter75_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter76_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter75_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter76_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter75_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter76_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter75_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter76_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter75_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter76_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter75_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter76_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter75_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter76_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter75_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter76_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter75_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter76_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter75_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter76_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter75_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter76_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter75_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter76_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter75_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter76_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter75_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter76_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter75_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter76_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter75_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter76_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter75_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter76_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter75_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter76_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter75_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter76_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter75_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter76_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter75_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter76_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter75_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter76_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter75_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter76_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter75_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter76_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter75_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter76_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter75_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter76_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter75_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter76_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter75_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter76_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter75_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter76_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter75_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter76_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter75_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter76_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter75_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter76_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter75_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter76_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter75_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter76_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter75_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter76_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter75_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter76_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter75_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter76_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter75_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter76_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter75_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter76_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter75_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter76_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter75_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter76_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter75_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter76_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter75_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter76_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter75_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter76_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter75_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter76_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter75_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter76_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter75_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter76_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter75_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter76_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter75_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter76_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter75_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter76_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter75_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter76_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter75_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter76_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter75_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter76_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter75_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter76_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter75_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter76_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter75_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter76_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter75_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter76_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter75_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter76_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter75_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter76_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter75_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter76_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter75_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter77_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter76_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter77_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter76_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter77_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter76_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter77_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter76_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter77_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter76_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter77_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter76_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter77_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter76_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter77_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter76_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter77_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter76_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter77_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter76_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter77_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter76_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter77_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter76_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter77_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter76_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter77_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter76_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter77_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter76_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter77_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter76_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter77_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter76_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter77_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter76_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter77_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter76_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter77_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter76_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter77_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter76_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter77_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter76_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter77_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter76_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter77_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter76_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter77_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter76_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter77_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter76_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter77_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter76_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter77_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter76_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter77_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter76_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter77_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter76_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter77_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter76_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter77_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter76_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter77_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter76_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter77_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter76_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter77_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter76_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter77_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter76_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter77_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter76_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter77_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter76_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter77_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter76_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter77_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter76_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter77_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter76_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter77_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter76_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter77_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter76_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter77_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter76_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter77_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter76_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter77_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter76_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter77_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter76_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter77_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter76_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter77_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter76_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter77_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter76_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter77_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter76_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter77_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter76_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter77_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter76_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter77_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter76_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter77_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter76_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter77_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter76_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter77_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter76_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter77_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter76_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter77_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter76_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter77_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter76_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter77_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter76_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter77_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter76_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter77_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter76_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter77_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter76_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter7_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter6_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter7_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter6_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter7_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter6_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter7_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter6_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter7_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter6_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter7_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter6_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter7_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter6_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter7_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter6_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter7_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter6_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter7_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter6_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter7_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter6_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter7_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter6_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter7_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter6_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter7_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter6_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter7_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter6_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter7_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter6_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter7_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter6_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter7_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter6_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter7_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter6_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter7_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter6_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter7_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter6_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter7_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter6_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter7_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter6_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter7_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter6_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter7_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter6_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter7_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter6_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter7_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter6_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter7_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter6_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter7_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter6_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter7_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter6_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter7_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter6_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter7_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter6_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter7_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter6_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter7_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter6_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter7_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter6_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter7_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter6_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter7_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter6_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter7_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter6_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter7_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter6_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter7_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter6_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter7_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter6_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter7_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter6_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter7_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter6_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter7_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter6_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter7_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter6_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter7_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter6_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter7_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter6_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter7_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter6_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter7_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter6_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter7_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter6_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter7_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter6_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter7_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter6_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter7_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter6_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter7_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter6_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter7_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter6_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter7_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter6_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter7_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter6_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter7_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter6_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter7_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter6_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter7_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter6_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter7_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter6_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter7_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter6_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter7_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter6_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter7_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter6_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter8_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter7_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter8_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter7_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter8_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter7_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter8_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter7_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter8_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter7_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter8_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter7_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter8_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter7_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter8_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter7_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter8_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter7_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter8_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter7_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter8_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter7_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter8_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter7_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter8_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter7_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter8_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter7_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter8_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter7_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter8_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter7_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter8_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter7_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter8_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter7_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter8_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter7_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter8_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter7_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter8_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter7_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter8_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter7_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter8_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter7_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter8_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter7_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter8_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter7_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter8_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter7_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter8_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter7_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter8_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter7_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter8_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter7_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter8_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter7_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter8_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter7_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter8_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter7_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter8_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter7_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter8_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter7_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter8_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter7_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter8_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter7_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter8_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter7_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter8_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter7_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter8_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter7_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter8_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter7_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter8_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter7_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter8_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter7_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter8_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter7_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter8_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter7_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter8_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter7_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter8_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter7_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter8_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter7_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter8_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter7_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter8_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter7_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter8_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter7_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter8_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter7_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter8_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter7_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter8_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter7_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter8_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter7_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter8_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter7_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter8_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter7_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter8_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter7_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter8_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter7_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter8_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter7_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter8_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter7_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter8_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter7_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter8_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter7_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter8_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter7_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter8_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter7_write_flag_0_reg_623;
            ap_phi_reg_pp0_iter9_phi_ln112_10_reg_1568 <= ap_phi_reg_pp0_iter8_phi_ln112_10_reg_1568;
            ap_phi_reg_pp0_iter9_phi_ln112_11_reg_1583 <= ap_phi_reg_pp0_iter8_phi_ln112_11_reg_1583;
            ap_phi_reg_pp0_iter9_phi_ln112_12_reg_1598 <= ap_phi_reg_pp0_iter8_phi_ln112_12_reg_1598;
            ap_phi_reg_pp0_iter9_phi_ln112_13_reg_1613 <= ap_phi_reg_pp0_iter8_phi_ln112_13_reg_1613;
            ap_phi_reg_pp0_iter9_phi_ln112_14_reg_1628 <= ap_phi_reg_pp0_iter8_phi_ln112_14_reg_1628;
            ap_phi_reg_pp0_iter9_phi_ln112_15_reg_1643 <= ap_phi_reg_pp0_iter8_phi_ln112_15_reg_1643;
            ap_phi_reg_pp0_iter9_phi_ln112_1_reg_1673 <= ap_phi_reg_pp0_iter8_phi_ln112_1_reg_1673;
            ap_phi_reg_pp0_iter9_phi_ln112_2_reg_1688 <= ap_phi_reg_pp0_iter8_phi_ln112_2_reg_1688;
            ap_phi_reg_pp0_iter9_phi_ln112_3_reg_1703 <= ap_phi_reg_pp0_iter8_phi_ln112_3_reg_1703;
            ap_phi_reg_pp0_iter9_phi_ln112_4_reg_1478 <= ap_phi_reg_pp0_iter8_phi_ln112_4_reg_1478;
            ap_phi_reg_pp0_iter9_phi_ln112_5_reg_1493 <= ap_phi_reg_pp0_iter8_phi_ln112_5_reg_1493;
            ap_phi_reg_pp0_iter9_phi_ln112_6_reg_1508 <= ap_phi_reg_pp0_iter8_phi_ln112_6_reg_1508;
            ap_phi_reg_pp0_iter9_phi_ln112_7_reg_1523 <= ap_phi_reg_pp0_iter8_phi_ln112_7_reg_1523;
            ap_phi_reg_pp0_iter9_phi_ln112_8_reg_1538 <= ap_phi_reg_pp0_iter8_phi_ln112_8_reg_1538;
            ap_phi_reg_pp0_iter9_phi_ln112_9_reg_1553 <= ap_phi_reg_pp0_iter8_phi_ln112_9_reg_1553;
            ap_phi_reg_pp0_iter9_phi_ln112_reg_1658 <= ap_phi_reg_pp0_iter8_phi_ln112_reg_1658;
            ap_phi_reg_pp0_iter9_write_flag101_0_reg_1212 <= ap_phi_reg_pp0_iter8_write_flag101_0_reg_1212;
            ap_phi_reg_pp0_iter9_write_flag104_0_reg_1193 <= ap_phi_reg_pp0_iter8_write_flag104_0_reg_1193;
            ap_phi_reg_pp0_iter9_write_flag107_0_reg_1174 <= ap_phi_reg_pp0_iter8_write_flag107_0_reg_1174;
            ap_phi_reg_pp0_iter9_write_flag110_0_reg_1307 <= ap_phi_reg_pp0_iter8_write_flag110_0_reg_1307;
            ap_phi_reg_pp0_iter9_write_flag113_0_reg_1288 <= ap_phi_reg_pp0_iter8_write_flag113_0_reg_1288;
            ap_phi_reg_pp0_iter9_write_flag116_0_reg_1269 <= ap_phi_reg_pp0_iter8_write_flag116_0_reg_1269;
            ap_phi_reg_pp0_iter9_write_flag119_0_reg_1250 <= ap_phi_reg_pp0_iter8_write_flag119_0_reg_1250;
            ap_phi_reg_pp0_iter9_write_flag11_0_reg_566 <= ap_phi_reg_pp0_iter8_write_flag11_0_reg_566;
            ap_phi_reg_pp0_iter9_write_flag122_0_reg_1383 <= ap_phi_reg_pp0_iter8_write_flag122_0_reg_1383;
            ap_phi_reg_pp0_iter9_write_flag125_0_reg_1345 <= ap_phi_reg_pp0_iter8_write_flag125_0_reg_1345;
            ap_phi_reg_pp0_iter9_write_flag128_0_reg_1326 <= ap_phi_reg_pp0_iter8_write_flag128_0_reg_1326;
            ap_phi_reg_pp0_iter9_write_flag131_0_reg_1364 <= ap_phi_reg_pp0_iter8_write_flag131_0_reg_1364;
            ap_phi_reg_pp0_iter9_write_flag134_0_reg_1402 <= ap_phi_reg_pp0_iter8_write_flag134_0_reg_1402;
            ap_phi_reg_pp0_iter9_write_flag137_0_reg_1421 <= ap_phi_reg_pp0_iter8_write_flag137_0_reg_1421;
            ap_phi_reg_pp0_iter9_write_flag140_0_reg_1440 <= ap_phi_reg_pp0_iter8_write_flag140_0_reg_1440;
            ap_phi_reg_pp0_iter9_write_flag143_0_reg_1459 <= ap_phi_reg_pp0_iter8_write_flag143_0_reg_1459;
            ap_phi_reg_pp0_iter9_write_flag14_0_reg_699 <= ap_phi_reg_pp0_iter8_write_flag14_0_reg_699;
            ap_phi_reg_pp0_iter9_write_flag17_0_reg_680 <= ap_phi_reg_pp0_iter8_write_flag17_0_reg_680;
            ap_phi_reg_pp0_iter9_write_flag20_0_reg_661 <= ap_phi_reg_pp0_iter8_write_flag20_0_reg_661;
            ap_phi_reg_pp0_iter9_write_flag23_0_reg_642 <= ap_phi_reg_pp0_iter8_write_flag23_0_reg_642;
            ap_phi_reg_pp0_iter9_write_flag26_0_reg_775 <= ap_phi_reg_pp0_iter8_write_flag26_0_reg_775;
            ap_phi_reg_pp0_iter9_write_flag29_0_reg_756 <= ap_phi_reg_pp0_iter8_write_flag29_0_reg_756;
            ap_phi_reg_pp0_iter9_write_flag32_0_reg_718 <= ap_phi_reg_pp0_iter8_write_flag32_0_reg_718;
            ap_phi_reg_pp0_iter9_write_flag35_0_reg_737 <= ap_phi_reg_pp0_iter8_write_flag35_0_reg_737;
            ap_phi_reg_pp0_iter9_write_flag38_0_reg_794 <= ap_phi_reg_pp0_iter8_write_flag38_0_reg_794;
            ap_phi_reg_pp0_iter9_write_flag41_0_reg_813 <= ap_phi_reg_pp0_iter8_write_flag41_0_reg_813;
            ap_phi_reg_pp0_iter9_write_flag44_0_reg_832 <= ap_phi_reg_pp0_iter8_write_flag44_0_reg_832;
            ap_phi_reg_pp0_iter9_write_flag47_0_reg_851 <= ap_phi_reg_pp0_iter8_write_flag47_0_reg_851;
            ap_phi_reg_pp0_iter9_write_flag4_0_reg_604 <= ap_phi_reg_pp0_iter8_write_flag4_0_reg_604;
            ap_phi_reg_pp0_iter9_write_flag50_0_reg_870 <= ap_phi_reg_pp0_iter8_write_flag50_0_reg_870;
            ap_phi_reg_pp0_iter9_write_flag53_0_reg_889 <= ap_phi_reg_pp0_iter8_write_flag53_0_reg_889;
            ap_phi_reg_pp0_iter9_write_flag56_0_reg_908 <= ap_phi_reg_pp0_iter8_write_flag56_0_reg_908;
            ap_phi_reg_pp0_iter9_write_flag59_0_reg_927 <= ap_phi_reg_pp0_iter8_write_flag59_0_reg_927;
            ap_phi_reg_pp0_iter9_write_flag62_0_reg_946 <= ap_phi_reg_pp0_iter8_write_flag62_0_reg_946;
            ap_phi_reg_pp0_iter9_write_flag65_0_reg_965 <= ap_phi_reg_pp0_iter8_write_flag65_0_reg_965;
            ap_phi_reg_pp0_iter9_write_flag68_0_reg_984 <= ap_phi_reg_pp0_iter8_write_flag68_0_reg_984;
            ap_phi_reg_pp0_iter9_write_flag71_0_reg_1003 <= ap_phi_reg_pp0_iter8_write_flag71_0_reg_1003;
            ap_phi_reg_pp0_iter9_write_flag74_0_reg_1022 <= ap_phi_reg_pp0_iter8_write_flag74_0_reg_1022;
            ap_phi_reg_pp0_iter9_write_flag77_0_reg_1041 <= ap_phi_reg_pp0_iter8_write_flag77_0_reg_1041;
            ap_phi_reg_pp0_iter9_write_flag80_0_reg_1060 <= ap_phi_reg_pp0_iter8_write_flag80_0_reg_1060;
            ap_phi_reg_pp0_iter9_write_flag83_0_reg_1079 <= ap_phi_reg_pp0_iter8_write_flag83_0_reg_1079;
            ap_phi_reg_pp0_iter9_write_flag86_0_reg_1098 <= ap_phi_reg_pp0_iter8_write_flag86_0_reg_1098;
            ap_phi_reg_pp0_iter9_write_flag89_0_reg_1117 <= ap_phi_reg_pp0_iter8_write_flag89_0_reg_1117;
            ap_phi_reg_pp0_iter9_write_flag8_0_reg_585 <= ap_phi_reg_pp0_iter8_write_flag8_0_reg_585;
            ap_phi_reg_pp0_iter9_write_flag92_0_reg_1136 <= ap_phi_reg_pp0_iter8_write_flag92_0_reg_1136;
            ap_phi_reg_pp0_iter9_write_flag95_0_reg_1155 <= ap_phi_reg_pp0_iter8_write_flag95_0_reg_1155;
            ap_phi_reg_pp0_iter9_write_flag98_0_reg_1231 <= ap_phi_reg_pp0_iter8_write_flag98_0_reg_1231;
            ap_phi_reg_pp0_iter9_write_flag_0_reg_623 <= ap_phi_reg_pp0_iter8_write_flag_0_reg_623;
            mul_i1_0_0_1_reg_3352 <= grp_fu_2107_p2;
            mul_i1_0_0_1_reg_3352_pp0_iter21_reg <= mul_i1_0_0_1_reg_3352;
            mul_i1_0_0_1_reg_3352_pp0_iter22_reg <= mul_i1_0_0_1_reg_3352_pp0_iter21_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter23_reg <= mul_i1_0_0_1_reg_3352_pp0_iter22_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter24_reg <= mul_i1_0_0_1_reg_3352_pp0_iter23_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter25_reg <= mul_i1_0_0_1_reg_3352_pp0_iter24_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter26_reg <= mul_i1_0_0_1_reg_3352_pp0_iter25_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter27_reg <= mul_i1_0_0_1_reg_3352_pp0_iter26_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter28_reg <= mul_i1_0_0_1_reg_3352_pp0_iter27_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter29_reg <= mul_i1_0_0_1_reg_3352_pp0_iter28_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter30_reg <= mul_i1_0_0_1_reg_3352_pp0_iter29_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter31_reg <= mul_i1_0_0_1_reg_3352_pp0_iter30_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter32_reg <= mul_i1_0_0_1_reg_3352_pp0_iter31_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter33_reg <= mul_i1_0_0_1_reg_3352_pp0_iter32_reg;
            mul_i1_0_0_1_reg_3352_pp0_iter34_reg <= mul_i1_0_0_1_reg_3352_pp0_iter33_reg;
            mul_i1_0_0_2_reg_3408 <= grp_fu_2132_p2;
            mul_i1_0_0_3_reg_3456 <= grp_fu_2147_p2;
            mul_i1_0_0_3_reg_3456_pp0_iter35_reg <= mul_i1_0_0_3_reg_3456;
            mul_i1_0_0_3_reg_3456_pp0_iter36_reg <= mul_i1_0_0_3_reg_3456_pp0_iter35_reg;
            mul_i1_0_0_3_reg_3456_pp0_iter37_reg <= mul_i1_0_0_3_reg_3456_pp0_iter36_reg;
            mul_i1_0_0_3_reg_3456_pp0_iter38_reg <= mul_i1_0_0_3_reg_3456_pp0_iter37_reg;
            mul_i1_0_0_3_reg_3456_pp0_iter39_reg <= mul_i1_0_0_3_reg_3456_pp0_iter38_reg;
            mul_i1_0_0_3_reg_3456_pp0_iter40_reg <= mul_i1_0_0_3_reg_3456_pp0_iter39_reg;
            mul_i1_0_0_3_reg_3456_pp0_iter41_reg <= mul_i1_0_0_3_reg_3456_pp0_iter40_reg;
            mul_i1_0_1_reg_3360 <= grp_fu_2112_p2;
            mul_i1_1_0_1_reg_3365 <= grp_fu_2117_p2;
            mul_i1_1_0_1_reg_3365_pp0_iter21_reg <= mul_i1_1_0_1_reg_3365;
            mul_i1_1_0_1_reg_3365_pp0_iter22_reg <= mul_i1_1_0_1_reg_3365_pp0_iter21_reg;
            mul_i1_1_0_1_reg_3365_pp0_iter23_reg <= mul_i1_1_0_1_reg_3365_pp0_iter22_reg;
            mul_i1_1_0_1_reg_3365_pp0_iter24_reg <= mul_i1_1_0_1_reg_3365_pp0_iter23_reg;
            mul_i1_1_0_1_reg_3365_pp0_iter25_reg <= mul_i1_1_0_1_reg_3365_pp0_iter24_reg;
            mul_i1_1_0_1_reg_3365_pp0_iter26_reg <= mul_i1_1_0_1_reg_3365_pp0_iter25_reg;
            mul_i1_1_0_1_reg_3365_pp0_iter27_reg <= mul_i1_1_0_1_reg_3365_pp0_iter26_reg;
            mul_i1_1_0_2_reg_3424 <= grp_fu_2137_p2;
            mul_i1_1_0_3_reg_3479 <= grp_fu_2152_p2;
            mul_i1_1_0_3_reg_3479_pp0_iter35_reg <= mul_i1_1_0_3_reg_3479;
            mul_i1_1_0_3_reg_3479_pp0_iter36_reg <= mul_i1_1_0_3_reg_3479_pp0_iter35_reg;
            mul_i1_1_0_3_reg_3479_pp0_iter37_reg <= mul_i1_1_0_3_reg_3479_pp0_iter36_reg;
            mul_i1_1_0_3_reg_3479_pp0_iter38_reg <= mul_i1_1_0_3_reg_3479_pp0_iter37_reg;
            mul_i1_1_0_3_reg_3479_pp0_iter39_reg <= mul_i1_1_0_3_reg_3479_pp0_iter38_reg;
            mul_i1_1_0_3_reg_3479_pp0_iter40_reg <= mul_i1_1_0_3_reg_3479_pp0_iter39_reg;
            mul_i1_1_0_3_reg_3479_pp0_iter41_reg <= mul_i1_1_0_3_reg_3479_pp0_iter40_reg;
            mul_i1_1_1_reg_3371 <= grp_fu_2122_p2;
            mul_i1_1_1_reg_3371_pp0_iter21_reg <= mul_i1_1_1_reg_3371;
            mul_i1_1_1_reg_3371_pp0_iter22_reg <= mul_i1_1_1_reg_3371_pp0_iter21_reg;
            mul_i1_1_1_reg_3371_pp0_iter23_reg <= mul_i1_1_1_reg_3371_pp0_iter22_reg;
            mul_i1_1_1_reg_3371_pp0_iter24_reg <= mul_i1_1_1_reg_3371_pp0_iter23_reg;
            mul_i1_1_1_reg_3371_pp0_iter25_reg <= mul_i1_1_1_reg_3371_pp0_iter24_reg;
            mul_i1_1_1_reg_3371_pp0_iter26_reg <= mul_i1_1_1_reg_3371_pp0_iter25_reg;
            mul_i1_1_1_reg_3371_pp0_iter27_reg <= mul_i1_1_1_reg_3371_pp0_iter26_reg;
            mul_i1_1_1_reg_3371_pp0_iter28_reg <= mul_i1_1_1_reg_3371_pp0_iter27_reg;
            mul_i1_1_1_reg_3371_pp0_iter29_reg <= mul_i1_1_1_reg_3371_pp0_iter28_reg;
            mul_i1_1_1_reg_3371_pp0_iter30_reg <= mul_i1_1_1_reg_3371_pp0_iter29_reg;
            mul_i1_1_1_reg_3371_pp0_iter31_reg <= mul_i1_1_1_reg_3371_pp0_iter30_reg;
            mul_i1_1_1_reg_3371_pp0_iter32_reg <= mul_i1_1_1_reg_3371_pp0_iter31_reg;
            mul_i1_1_1_reg_3371_pp0_iter33_reg <= mul_i1_1_1_reg_3371_pp0_iter32_reg;
            mul_i1_1_1_reg_3371_pp0_iter34_reg <= mul_i1_1_1_reg_3371_pp0_iter33_reg;
            mul_i1_2_0_1_reg_3378 <= grp_fu_2127_p2;
            mul_i1_2_0_1_reg_3378_pp0_iter21_reg <= mul_i1_2_0_1_reg_3378;
            mul_i1_2_0_1_reg_3378_pp0_iter22_reg <= mul_i1_2_0_1_reg_3378_pp0_iter21_reg;
            mul_i1_2_0_1_reg_3378_pp0_iter23_reg <= mul_i1_2_0_1_reg_3378_pp0_iter22_reg;
            mul_i1_2_0_1_reg_3378_pp0_iter24_reg <= mul_i1_2_0_1_reg_3378_pp0_iter23_reg;
            mul_i1_2_0_1_reg_3378_pp0_iter25_reg <= mul_i1_2_0_1_reg_3378_pp0_iter24_reg;
            mul_i1_2_0_1_reg_3378_pp0_iter26_reg <= mul_i1_2_0_1_reg_3378_pp0_iter25_reg;
            mul_i1_2_0_1_reg_3378_pp0_iter27_reg <= mul_i1_2_0_1_reg_3378_pp0_iter26_reg;
            mul_i1_2_0_2_reg_3440 <= grp_fu_2142_p2;
            mul_i1_2_0_3_reg_3502 <= grp_fu_2157_p2;
            mul_i1_2_0_3_reg_3502_pp0_iter35_reg <= mul_i1_2_0_3_reg_3502;
            mul_i1_2_0_3_reg_3502_pp0_iter36_reg <= mul_i1_2_0_3_reg_3502_pp0_iter35_reg;
            mul_i1_2_0_3_reg_3502_pp0_iter37_reg <= mul_i1_2_0_3_reg_3502_pp0_iter36_reg;
            mul_i1_2_0_3_reg_3502_pp0_iter38_reg <= mul_i1_2_0_3_reg_3502_pp0_iter37_reg;
            mul_i1_2_0_3_reg_3502_pp0_iter39_reg <= mul_i1_2_0_3_reg_3502_pp0_iter38_reg;
            mul_i1_2_0_3_reg_3502_pp0_iter40_reg <= mul_i1_2_0_3_reg_3502_pp0_iter39_reg;
            mul_i1_2_0_3_reg_3502_pp0_iter41_reg <= mul_i1_2_0_3_reg_3502_pp0_iter40_reg;
            mul_i1_2_1_2_reg_3514 <= grp_fu_2162_p2;
            mul_i2_0_0_1_reg_3666 <= grp_fu_2182_p2;
            mul_i2_0_0_2_reg_3735 <= grp_fu_2212_p2;
            mul_i2_0_0_3_reg_3816 <= grp_fu_2227_p2;
            mul_i2_0_1_reg_3646 <= grp_fu_2167_p2;
            mul_i2_0_2_1_reg_3679 <= grp_fu_2187_p2;
            mul_i2_1_0_1_reg_3689 <= grp_fu_2192_p2;
            mul_i2_1_0_2_reg_3762 <= grp_fu_2217_p2;
            mul_i2_1_0_3_reg_3843 <= grp_fu_2232_p2;
            mul_i2_1_1_reg_3651 <= grp_fu_2172_p2;
            mul_i2_1_2_1_reg_3702 <= grp_fu_2197_p2;
            mul_i2_2_0_1_reg_3712 <= grp_fu_2202_p2;
            mul_i2_2_0_2_reg_3789 <= grp_fu_2222_p2;
            mul_i2_2_0_3_reg_3870 <= grp_fu_2237_p2;
            mul_i2_2_1_reg_3656 <= grp_fu_2177_p2;
            mul_i2_2_2_1_reg_3725 <= grp_fu_2207_p2;
            mul_i_0_0_3_reg_3287 <= grp_fu_2089_p2;
            mul_i_1_0_3_reg_3293 <= grp_fu_2095_p2;
            mul_i_2_0_3_reg_3299 <= grp_fu_2101_p2;
            mul_i_2_0_3_reg_3299_pp0_iter10_reg <= mul_i_2_0_3_reg_3299_pp0_iter9_reg;
            mul_i_2_0_3_reg_3299_pp0_iter11_reg <= mul_i_2_0_3_reg_3299_pp0_iter10_reg;
            mul_i_2_0_3_reg_3299_pp0_iter12_reg <= mul_i_2_0_3_reg_3299_pp0_iter11_reg;
            mul_i_2_0_3_reg_3299_pp0_iter13_reg <= mul_i_2_0_3_reg_3299_pp0_iter12_reg;
            mul_i_2_0_3_reg_3299_pp0_iter7_reg <= mul_i_2_0_3_reg_3299;
            mul_i_2_0_3_reg_3299_pp0_iter8_reg <= mul_i_2_0_3_reg_3299_pp0_iter7_reg;
            mul_i_2_0_3_reg_3299_pp0_iter9_reg <= mul_i_2_0_3_reg_3299_pp0_iter8_reg;
            p_read64_reg_3264 <= p_read_int_reg;
            p_read64_reg_3264_pp0_iter10_reg <= p_read64_reg_3264_pp0_iter9_reg;
            p_read64_reg_3264_pp0_iter11_reg <= p_read64_reg_3264_pp0_iter10_reg;
            p_read64_reg_3264_pp0_iter12_reg <= p_read64_reg_3264_pp0_iter11_reg;
            p_read64_reg_3264_pp0_iter13_reg <= p_read64_reg_3264_pp0_iter12_reg;
            p_read64_reg_3264_pp0_iter14_reg <= p_read64_reg_3264_pp0_iter13_reg;
            p_read64_reg_3264_pp0_iter15_reg <= p_read64_reg_3264_pp0_iter14_reg;
            p_read64_reg_3264_pp0_iter16_reg <= p_read64_reg_3264_pp0_iter15_reg;
            p_read64_reg_3264_pp0_iter17_reg <= p_read64_reg_3264_pp0_iter16_reg;
            p_read64_reg_3264_pp0_iter18_reg <= p_read64_reg_3264_pp0_iter17_reg;
            p_read64_reg_3264_pp0_iter19_reg <= p_read64_reg_3264_pp0_iter18_reg;
            p_read64_reg_3264_pp0_iter1_reg <= p_read64_reg_3264;
            p_read64_reg_3264_pp0_iter20_reg <= p_read64_reg_3264_pp0_iter19_reg;
            p_read64_reg_3264_pp0_iter21_reg <= p_read64_reg_3264_pp0_iter20_reg;
            p_read64_reg_3264_pp0_iter22_reg <= p_read64_reg_3264_pp0_iter21_reg;
            p_read64_reg_3264_pp0_iter23_reg <= p_read64_reg_3264_pp0_iter22_reg;
            p_read64_reg_3264_pp0_iter24_reg <= p_read64_reg_3264_pp0_iter23_reg;
            p_read64_reg_3264_pp0_iter25_reg <= p_read64_reg_3264_pp0_iter24_reg;
            p_read64_reg_3264_pp0_iter26_reg <= p_read64_reg_3264_pp0_iter25_reg;
            p_read64_reg_3264_pp0_iter27_reg <= p_read64_reg_3264_pp0_iter26_reg;
            p_read64_reg_3264_pp0_iter28_reg <= p_read64_reg_3264_pp0_iter27_reg;
            p_read64_reg_3264_pp0_iter29_reg <= p_read64_reg_3264_pp0_iter28_reg;
            p_read64_reg_3264_pp0_iter2_reg <= p_read64_reg_3264_pp0_iter1_reg;
            p_read64_reg_3264_pp0_iter30_reg <= p_read64_reg_3264_pp0_iter29_reg;
            p_read64_reg_3264_pp0_iter31_reg <= p_read64_reg_3264_pp0_iter30_reg;
            p_read64_reg_3264_pp0_iter32_reg <= p_read64_reg_3264_pp0_iter31_reg;
            p_read64_reg_3264_pp0_iter33_reg <= p_read64_reg_3264_pp0_iter32_reg;
            p_read64_reg_3264_pp0_iter34_reg <= p_read64_reg_3264_pp0_iter33_reg;
            p_read64_reg_3264_pp0_iter35_reg <= p_read64_reg_3264_pp0_iter34_reg;
            p_read64_reg_3264_pp0_iter36_reg <= p_read64_reg_3264_pp0_iter35_reg;
            p_read64_reg_3264_pp0_iter37_reg <= p_read64_reg_3264_pp0_iter36_reg;
            p_read64_reg_3264_pp0_iter38_reg <= p_read64_reg_3264_pp0_iter37_reg;
            p_read64_reg_3264_pp0_iter39_reg <= p_read64_reg_3264_pp0_iter38_reg;
            p_read64_reg_3264_pp0_iter3_reg <= p_read64_reg_3264_pp0_iter2_reg;
            p_read64_reg_3264_pp0_iter40_reg <= p_read64_reg_3264_pp0_iter39_reg;
            p_read64_reg_3264_pp0_iter41_reg <= p_read64_reg_3264_pp0_iter40_reg;
            p_read64_reg_3264_pp0_iter42_reg <= p_read64_reg_3264_pp0_iter41_reg;
            p_read64_reg_3264_pp0_iter43_reg <= p_read64_reg_3264_pp0_iter42_reg;
            p_read64_reg_3264_pp0_iter44_reg <= p_read64_reg_3264_pp0_iter43_reg;
            p_read64_reg_3264_pp0_iter45_reg <= p_read64_reg_3264_pp0_iter44_reg;
            p_read64_reg_3264_pp0_iter46_reg <= p_read64_reg_3264_pp0_iter45_reg;
            p_read64_reg_3264_pp0_iter47_reg <= p_read64_reg_3264_pp0_iter46_reg;
            p_read64_reg_3264_pp0_iter48_reg <= p_read64_reg_3264_pp0_iter47_reg;
            p_read64_reg_3264_pp0_iter49_reg <= p_read64_reg_3264_pp0_iter48_reg;
            p_read64_reg_3264_pp0_iter4_reg <= p_read64_reg_3264_pp0_iter3_reg;
            p_read64_reg_3264_pp0_iter50_reg <= p_read64_reg_3264_pp0_iter49_reg;
            p_read64_reg_3264_pp0_iter51_reg <= p_read64_reg_3264_pp0_iter50_reg;
            p_read64_reg_3264_pp0_iter52_reg <= p_read64_reg_3264_pp0_iter51_reg;
            p_read64_reg_3264_pp0_iter53_reg <= p_read64_reg_3264_pp0_iter52_reg;
            p_read64_reg_3264_pp0_iter54_reg <= p_read64_reg_3264_pp0_iter53_reg;
            p_read64_reg_3264_pp0_iter55_reg <= p_read64_reg_3264_pp0_iter54_reg;
            p_read64_reg_3264_pp0_iter56_reg <= p_read64_reg_3264_pp0_iter55_reg;
            p_read64_reg_3264_pp0_iter57_reg <= p_read64_reg_3264_pp0_iter56_reg;
            p_read64_reg_3264_pp0_iter58_reg <= p_read64_reg_3264_pp0_iter57_reg;
            p_read64_reg_3264_pp0_iter59_reg <= p_read64_reg_3264_pp0_iter58_reg;
            p_read64_reg_3264_pp0_iter5_reg <= p_read64_reg_3264_pp0_iter4_reg;
            p_read64_reg_3264_pp0_iter60_reg <= p_read64_reg_3264_pp0_iter59_reg;
            p_read64_reg_3264_pp0_iter61_reg <= p_read64_reg_3264_pp0_iter60_reg;
            p_read64_reg_3264_pp0_iter62_reg <= p_read64_reg_3264_pp0_iter61_reg;
            p_read64_reg_3264_pp0_iter63_reg <= p_read64_reg_3264_pp0_iter62_reg;
            p_read64_reg_3264_pp0_iter64_reg <= p_read64_reg_3264_pp0_iter63_reg;
            p_read64_reg_3264_pp0_iter65_reg <= p_read64_reg_3264_pp0_iter64_reg;
            p_read64_reg_3264_pp0_iter66_reg <= p_read64_reg_3264_pp0_iter65_reg;
            p_read64_reg_3264_pp0_iter67_reg <= p_read64_reg_3264_pp0_iter66_reg;
            p_read64_reg_3264_pp0_iter68_reg <= p_read64_reg_3264_pp0_iter67_reg;
            p_read64_reg_3264_pp0_iter69_reg <= p_read64_reg_3264_pp0_iter68_reg;
            p_read64_reg_3264_pp0_iter6_reg <= p_read64_reg_3264_pp0_iter5_reg;
            p_read64_reg_3264_pp0_iter70_reg <= p_read64_reg_3264_pp0_iter69_reg;
            p_read64_reg_3264_pp0_iter71_reg <= p_read64_reg_3264_pp0_iter70_reg;
            p_read64_reg_3264_pp0_iter72_reg <= p_read64_reg_3264_pp0_iter71_reg;
            p_read64_reg_3264_pp0_iter73_reg <= p_read64_reg_3264_pp0_iter72_reg;
            p_read64_reg_3264_pp0_iter74_reg <= p_read64_reg_3264_pp0_iter73_reg;
            p_read64_reg_3264_pp0_iter75_reg <= p_read64_reg_3264_pp0_iter74_reg;
            p_read64_reg_3264_pp0_iter76_reg <= p_read64_reg_3264_pp0_iter75_reg;
            p_read64_reg_3264_pp0_iter7_reg <= p_read64_reg_3264_pp0_iter6_reg;
            p_read64_reg_3264_pp0_iter8_reg <= p_read64_reg_3264_pp0_iter7_reg;
            p_read64_reg_3264_pp0_iter9_reg <= p_read64_reg_3264_pp0_iter8_reg;
            p_read_17_reg_3029 <= p_read47_int_reg;
            p_read_17_reg_3029_pp0_iter10_reg <= p_read_17_reg_3029_pp0_iter9_reg;
            p_read_17_reg_3029_pp0_iter11_reg <= p_read_17_reg_3029_pp0_iter10_reg;
            p_read_17_reg_3029_pp0_iter12_reg <= p_read_17_reg_3029_pp0_iter11_reg;
            p_read_17_reg_3029_pp0_iter13_reg <= p_read_17_reg_3029_pp0_iter12_reg;
            p_read_17_reg_3029_pp0_iter14_reg <= p_read_17_reg_3029_pp0_iter13_reg;
            p_read_17_reg_3029_pp0_iter15_reg <= p_read_17_reg_3029_pp0_iter14_reg;
            p_read_17_reg_3029_pp0_iter16_reg <= p_read_17_reg_3029_pp0_iter15_reg;
            p_read_17_reg_3029_pp0_iter17_reg <= p_read_17_reg_3029_pp0_iter16_reg;
            p_read_17_reg_3029_pp0_iter18_reg <= p_read_17_reg_3029_pp0_iter17_reg;
            p_read_17_reg_3029_pp0_iter19_reg <= p_read_17_reg_3029_pp0_iter18_reg;
            p_read_17_reg_3029_pp0_iter1_reg <= p_read_17_reg_3029;
            p_read_17_reg_3029_pp0_iter20_reg <= p_read_17_reg_3029_pp0_iter19_reg;
            p_read_17_reg_3029_pp0_iter21_reg <= p_read_17_reg_3029_pp0_iter20_reg;
            p_read_17_reg_3029_pp0_iter22_reg <= p_read_17_reg_3029_pp0_iter21_reg;
            p_read_17_reg_3029_pp0_iter23_reg <= p_read_17_reg_3029_pp0_iter22_reg;
            p_read_17_reg_3029_pp0_iter24_reg <= p_read_17_reg_3029_pp0_iter23_reg;
            p_read_17_reg_3029_pp0_iter25_reg <= p_read_17_reg_3029_pp0_iter24_reg;
            p_read_17_reg_3029_pp0_iter26_reg <= p_read_17_reg_3029_pp0_iter25_reg;
            p_read_17_reg_3029_pp0_iter27_reg <= p_read_17_reg_3029_pp0_iter26_reg;
            p_read_17_reg_3029_pp0_iter28_reg <= p_read_17_reg_3029_pp0_iter27_reg;
            p_read_17_reg_3029_pp0_iter29_reg <= p_read_17_reg_3029_pp0_iter28_reg;
            p_read_17_reg_3029_pp0_iter2_reg <= p_read_17_reg_3029_pp0_iter1_reg;
            p_read_17_reg_3029_pp0_iter30_reg <= p_read_17_reg_3029_pp0_iter29_reg;
            p_read_17_reg_3029_pp0_iter31_reg <= p_read_17_reg_3029_pp0_iter30_reg;
            p_read_17_reg_3029_pp0_iter32_reg <= p_read_17_reg_3029_pp0_iter31_reg;
            p_read_17_reg_3029_pp0_iter33_reg <= p_read_17_reg_3029_pp0_iter32_reg;
            p_read_17_reg_3029_pp0_iter34_reg <= p_read_17_reg_3029_pp0_iter33_reg;
            p_read_17_reg_3029_pp0_iter35_reg <= p_read_17_reg_3029_pp0_iter34_reg;
            p_read_17_reg_3029_pp0_iter36_reg <= p_read_17_reg_3029_pp0_iter35_reg;
            p_read_17_reg_3029_pp0_iter37_reg <= p_read_17_reg_3029_pp0_iter36_reg;
            p_read_17_reg_3029_pp0_iter38_reg <= p_read_17_reg_3029_pp0_iter37_reg;
            p_read_17_reg_3029_pp0_iter39_reg <= p_read_17_reg_3029_pp0_iter38_reg;
            p_read_17_reg_3029_pp0_iter3_reg <= p_read_17_reg_3029_pp0_iter2_reg;
            p_read_17_reg_3029_pp0_iter40_reg <= p_read_17_reg_3029_pp0_iter39_reg;
            p_read_17_reg_3029_pp0_iter41_reg <= p_read_17_reg_3029_pp0_iter40_reg;
            p_read_17_reg_3029_pp0_iter42_reg <= p_read_17_reg_3029_pp0_iter41_reg;
            p_read_17_reg_3029_pp0_iter43_reg <= p_read_17_reg_3029_pp0_iter42_reg;
            p_read_17_reg_3029_pp0_iter44_reg <= p_read_17_reg_3029_pp0_iter43_reg;
            p_read_17_reg_3029_pp0_iter45_reg <= p_read_17_reg_3029_pp0_iter44_reg;
            p_read_17_reg_3029_pp0_iter46_reg <= p_read_17_reg_3029_pp0_iter45_reg;
            p_read_17_reg_3029_pp0_iter47_reg <= p_read_17_reg_3029_pp0_iter46_reg;
            p_read_17_reg_3029_pp0_iter48_reg <= p_read_17_reg_3029_pp0_iter47_reg;
            p_read_17_reg_3029_pp0_iter49_reg <= p_read_17_reg_3029_pp0_iter48_reg;
            p_read_17_reg_3029_pp0_iter4_reg <= p_read_17_reg_3029_pp0_iter3_reg;
            p_read_17_reg_3029_pp0_iter50_reg <= p_read_17_reg_3029_pp0_iter49_reg;
            p_read_17_reg_3029_pp0_iter51_reg <= p_read_17_reg_3029_pp0_iter50_reg;
            p_read_17_reg_3029_pp0_iter52_reg <= p_read_17_reg_3029_pp0_iter51_reg;
            p_read_17_reg_3029_pp0_iter53_reg <= p_read_17_reg_3029_pp0_iter52_reg;
            p_read_17_reg_3029_pp0_iter54_reg <= p_read_17_reg_3029_pp0_iter53_reg;
            p_read_17_reg_3029_pp0_iter55_reg <= p_read_17_reg_3029_pp0_iter54_reg;
            p_read_17_reg_3029_pp0_iter56_reg <= p_read_17_reg_3029_pp0_iter55_reg;
            p_read_17_reg_3029_pp0_iter57_reg <= p_read_17_reg_3029_pp0_iter56_reg;
            p_read_17_reg_3029_pp0_iter58_reg <= p_read_17_reg_3029_pp0_iter57_reg;
            p_read_17_reg_3029_pp0_iter59_reg <= p_read_17_reg_3029_pp0_iter58_reg;
            p_read_17_reg_3029_pp0_iter5_reg <= p_read_17_reg_3029_pp0_iter4_reg;
            p_read_17_reg_3029_pp0_iter60_reg <= p_read_17_reg_3029_pp0_iter59_reg;
            p_read_17_reg_3029_pp0_iter61_reg <= p_read_17_reg_3029_pp0_iter60_reg;
            p_read_17_reg_3029_pp0_iter62_reg <= p_read_17_reg_3029_pp0_iter61_reg;
            p_read_17_reg_3029_pp0_iter63_reg <= p_read_17_reg_3029_pp0_iter62_reg;
            p_read_17_reg_3029_pp0_iter64_reg <= p_read_17_reg_3029_pp0_iter63_reg;
            p_read_17_reg_3029_pp0_iter65_reg <= p_read_17_reg_3029_pp0_iter64_reg;
            p_read_17_reg_3029_pp0_iter66_reg <= p_read_17_reg_3029_pp0_iter65_reg;
            p_read_17_reg_3029_pp0_iter67_reg <= p_read_17_reg_3029_pp0_iter66_reg;
            p_read_17_reg_3029_pp0_iter68_reg <= p_read_17_reg_3029_pp0_iter67_reg;
            p_read_17_reg_3029_pp0_iter69_reg <= p_read_17_reg_3029_pp0_iter68_reg;
            p_read_17_reg_3029_pp0_iter6_reg <= p_read_17_reg_3029_pp0_iter5_reg;
            p_read_17_reg_3029_pp0_iter70_reg <= p_read_17_reg_3029_pp0_iter69_reg;
            p_read_17_reg_3029_pp0_iter71_reg <= p_read_17_reg_3029_pp0_iter70_reg;
            p_read_17_reg_3029_pp0_iter72_reg <= p_read_17_reg_3029_pp0_iter71_reg;
            p_read_17_reg_3029_pp0_iter73_reg <= p_read_17_reg_3029_pp0_iter72_reg;
            p_read_17_reg_3029_pp0_iter74_reg <= p_read_17_reg_3029_pp0_iter73_reg;
            p_read_17_reg_3029_pp0_iter75_reg <= p_read_17_reg_3029_pp0_iter74_reg;
            p_read_17_reg_3029_pp0_iter76_reg <= p_read_17_reg_3029_pp0_iter75_reg;
            p_read_17_reg_3029_pp0_iter7_reg <= p_read_17_reg_3029_pp0_iter6_reg;
            p_read_17_reg_3029_pp0_iter8_reg <= p_read_17_reg_3029_pp0_iter7_reg;
            p_read_17_reg_3029_pp0_iter9_reg <= p_read_17_reg_3029_pp0_iter8_reg;
            p_read_18_reg_3034 <= p_read46_int_reg;
            p_read_18_reg_3034_pp0_iter10_reg <= p_read_18_reg_3034_pp0_iter9_reg;
            p_read_18_reg_3034_pp0_iter11_reg <= p_read_18_reg_3034_pp0_iter10_reg;
            p_read_18_reg_3034_pp0_iter12_reg <= p_read_18_reg_3034_pp0_iter11_reg;
            p_read_18_reg_3034_pp0_iter13_reg <= p_read_18_reg_3034_pp0_iter12_reg;
            p_read_18_reg_3034_pp0_iter14_reg <= p_read_18_reg_3034_pp0_iter13_reg;
            p_read_18_reg_3034_pp0_iter15_reg <= p_read_18_reg_3034_pp0_iter14_reg;
            p_read_18_reg_3034_pp0_iter16_reg <= p_read_18_reg_3034_pp0_iter15_reg;
            p_read_18_reg_3034_pp0_iter17_reg <= p_read_18_reg_3034_pp0_iter16_reg;
            p_read_18_reg_3034_pp0_iter18_reg <= p_read_18_reg_3034_pp0_iter17_reg;
            p_read_18_reg_3034_pp0_iter19_reg <= p_read_18_reg_3034_pp0_iter18_reg;
            p_read_18_reg_3034_pp0_iter1_reg <= p_read_18_reg_3034;
            p_read_18_reg_3034_pp0_iter20_reg <= p_read_18_reg_3034_pp0_iter19_reg;
            p_read_18_reg_3034_pp0_iter21_reg <= p_read_18_reg_3034_pp0_iter20_reg;
            p_read_18_reg_3034_pp0_iter22_reg <= p_read_18_reg_3034_pp0_iter21_reg;
            p_read_18_reg_3034_pp0_iter23_reg <= p_read_18_reg_3034_pp0_iter22_reg;
            p_read_18_reg_3034_pp0_iter24_reg <= p_read_18_reg_3034_pp0_iter23_reg;
            p_read_18_reg_3034_pp0_iter25_reg <= p_read_18_reg_3034_pp0_iter24_reg;
            p_read_18_reg_3034_pp0_iter26_reg <= p_read_18_reg_3034_pp0_iter25_reg;
            p_read_18_reg_3034_pp0_iter27_reg <= p_read_18_reg_3034_pp0_iter26_reg;
            p_read_18_reg_3034_pp0_iter28_reg <= p_read_18_reg_3034_pp0_iter27_reg;
            p_read_18_reg_3034_pp0_iter29_reg <= p_read_18_reg_3034_pp0_iter28_reg;
            p_read_18_reg_3034_pp0_iter2_reg <= p_read_18_reg_3034_pp0_iter1_reg;
            p_read_18_reg_3034_pp0_iter30_reg <= p_read_18_reg_3034_pp0_iter29_reg;
            p_read_18_reg_3034_pp0_iter31_reg <= p_read_18_reg_3034_pp0_iter30_reg;
            p_read_18_reg_3034_pp0_iter32_reg <= p_read_18_reg_3034_pp0_iter31_reg;
            p_read_18_reg_3034_pp0_iter33_reg <= p_read_18_reg_3034_pp0_iter32_reg;
            p_read_18_reg_3034_pp0_iter34_reg <= p_read_18_reg_3034_pp0_iter33_reg;
            p_read_18_reg_3034_pp0_iter35_reg <= p_read_18_reg_3034_pp0_iter34_reg;
            p_read_18_reg_3034_pp0_iter36_reg <= p_read_18_reg_3034_pp0_iter35_reg;
            p_read_18_reg_3034_pp0_iter37_reg <= p_read_18_reg_3034_pp0_iter36_reg;
            p_read_18_reg_3034_pp0_iter38_reg <= p_read_18_reg_3034_pp0_iter37_reg;
            p_read_18_reg_3034_pp0_iter39_reg <= p_read_18_reg_3034_pp0_iter38_reg;
            p_read_18_reg_3034_pp0_iter3_reg <= p_read_18_reg_3034_pp0_iter2_reg;
            p_read_18_reg_3034_pp0_iter40_reg <= p_read_18_reg_3034_pp0_iter39_reg;
            p_read_18_reg_3034_pp0_iter41_reg <= p_read_18_reg_3034_pp0_iter40_reg;
            p_read_18_reg_3034_pp0_iter42_reg <= p_read_18_reg_3034_pp0_iter41_reg;
            p_read_18_reg_3034_pp0_iter43_reg <= p_read_18_reg_3034_pp0_iter42_reg;
            p_read_18_reg_3034_pp0_iter44_reg <= p_read_18_reg_3034_pp0_iter43_reg;
            p_read_18_reg_3034_pp0_iter45_reg <= p_read_18_reg_3034_pp0_iter44_reg;
            p_read_18_reg_3034_pp0_iter46_reg <= p_read_18_reg_3034_pp0_iter45_reg;
            p_read_18_reg_3034_pp0_iter47_reg <= p_read_18_reg_3034_pp0_iter46_reg;
            p_read_18_reg_3034_pp0_iter48_reg <= p_read_18_reg_3034_pp0_iter47_reg;
            p_read_18_reg_3034_pp0_iter49_reg <= p_read_18_reg_3034_pp0_iter48_reg;
            p_read_18_reg_3034_pp0_iter4_reg <= p_read_18_reg_3034_pp0_iter3_reg;
            p_read_18_reg_3034_pp0_iter50_reg <= p_read_18_reg_3034_pp0_iter49_reg;
            p_read_18_reg_3034_pp0_iter51_reg <= p_read_18_reg_3034_pp0_iter50_reg;
            p_read_18_reg_3034_pp0_iter52_reg <= p_read_18_reg_3034_pp0_iter51_reg;
            p_read_18_reg_3034_pp0_iter53_reg <= p_read_18_reg_3034_pp0_iter52_reg;
            p_read_18_reg_3034_pp0_iter54_reg <= p_read_18_reg_3034_pp0_iter53_reg;
            p_read_18_reg_3034_pp0_iter55_reg <= p_read_18_reg_3034_pp0_iter54_reg;
            p_read_18_reg_3034_pp0_iter56_reg <= p_read_18_reg_3034_pp0_iter55_reg;
            p_read_18_reg_3034_pp0_iter57_reg <= p_read_18_reg_3034_pp0_iter56_reg;
            p_read_18_reg_3034_pp0_iter58_reg <= p_read_18_reg_3034_pp0_iter57_reg;
            p_read_18_reg_3034_pp0_iter59_reg <= p_read_18_reg_3034_pp0_iter58_reg;
            p_read_18_reg_3034_pp0_iter5_reg <= p_read_18_reg_3034_pp0_iter4_reg;
            p_read_18_reg_3034_pp0_iter60_reg <= p_read_18_reg_3034_pp0_iter59_reg;
            p_read_18_reg_3034_pp0_iter61_reg <= p_read_18_reg_3034_pp0_iter60_reg;
            p_read_18_reg_3034_pp0_iter62_reg <= p_read_18_reg_3034_pp0_iter61_reg;
            p_read_18_reg_3034_pp0_iter63_reg <= p_read_18_reg_3034_pp0_iter62_reg;
            p_read_18_reg_3034_pp0_iter64_reg <= p_read_18_reg_3034_pp0_iter63_reg;
            p_read_18_reg_3034_pp0_iter65_reg <= p_read_18_reg_3034_pp0_iter64_reg;
            p_read_18_reg_3034_pp0_iter66_reg <= p_read_18_reg_3034_pp0_iter65_reg;
            p_read_18_reg_3034_pp0_iter67_reg <= p_read_18_reg_3034_pp0_iter66_reg;
            p_read_18_reg_3034_pp0_iter68_reg <= p_read_18_reg_3034_pp0_iter67_reg;
            p_read_18_reg_3034_pp0_iter69_reg <= p_read_18_reg_3034_pp0_iter68_reg;
            p_read_18_reg_3034_pp0_iter6_reg <= p_read_18_reg_3034_pp0_iter5_reg;
            p_read_18_reg_3034_pp0_iter70_reg <= p_read_18_reg_3034_pp0_iter69_reg;
            p_read_18_reg_3034_pp0_iter71_reg <= p_read_18_reg_3034_pp0_iter70_reg;
            p_read_18_reg_3034_pp0_iter72_reg <= p_read_18_reg_3034_pp0_iter71_reg;
            p_read_18_reg_3034_pp0_iter73_reg <= p_read_18_reg_3034_pp0_iter72_reg;
            p_read_18_reg_3034_pp0_iter74_reg <= p_read_18_reg_3034_pp0_iter73_reg;
            p_read_18_reg_3034_pp0_iter75_reg <= p_read_18_reg_3034_pp0_iter74_reg;
            p_read_18_reg_3034_pp0_iter76_reg <= p_read_18_reg_3034_pp0_iter75_reg;
            p_read_18_reg_3034_pp0_iter7_reg <= p_read_18_reg_3034_pp0_iter6_reg;
            p_read_18_reg_3034_pp0_iter8_reg <= p_read_18_reg_3034_pp0_iter7_reg;
            p_read_18_reg_3034_pp0_iter9_reg <= p_read_18_reg_3034_pp0_iter8_reg;
            p_read_19_reg_3039 <= p_read45_int_reg;
            p_read_19_reg_3039_pp0_iter10_reg <= p_read_19_reg_3039_pp0_iter9_reg;
            p_read_19_reg_3039_pp0_iter11_reg <= p_read_19_reg_3039_pp0_iter10_reg;
            p_read_19_reg_3039_pp0_iter12_reg <= p_read_19_reg_3039_pp0_iter11_reg;
            p_read_19_reg_3039_pp0_iter13_reg <= p_read_19_reg_3039_pp0_iter12_reg;
            p_read_19_reg_3039_pp0_iter14_reg <= p_read_19_reg_3039_pp0_iter13_reg;
            p_read_19_reg_3039_pp0_iter15_reg <= p_read_19_reg_3039_pp0_iter14_reg;
            p_read_19_reg_3039_pp0_iter16_reg <= p_read_19_reg_3039_pp0_iter15_reg;
            p_read_19_reg_3039_pp0_iter17_reg <= p_read_19_reg_3039_pp0_iter16_reg;
            p_read_19_reg_3039_pp0_iter18_reg <= p_read_19_reg_3039_pp0_iter17_reg;
            p_read_19_reg_3039_pp0_iter19_reg <= p_read_19_reg_3039_pp0_iter18_reg;
            p_read_19_reg_3039_pp0_iter1_reg <= p_read_19_reg_3039;
            p_read_19_reg_3039_pp0_iter20_reg <= p_read_19_reg_3039_pp0_iter19_reg;
            p_read_19_reg_3039_pp0_iter21_reg <= p_read_19_reg_3039_pp0_iter20_reg;
            p_read_19_reg_3039_pp0_iter22_reg <= p_read_19_reg_3039_pp0_iter21_reg;
            p_read_19_reg_3039_pp0_iter23_reg <= p_read_19_reg_3039_pp0_iter22_reg;
            p_read_19_reg_3039_pp0_iter24_reg <= p_read_19_reg_3039_pp0_iter23_reg;
            p_read_19_reg_3039_pp0_iter25_reg <= p_read_19_reg_3039_pp0_iter24_reg;
            p_read_19_reg_3039_pp0_iter26_reg <= p_read_19_reg_3039_pp0_iter25_reg;
            p_read_19_reg_3039_pp0_iter27_reg <= p_read_19_reg_3039_pp0_iter26_reg;
            p_read_19_reg_3039_pp0_iter28_reg <= p_read_19_reg_3039_pp0_iter27_reg;
            p_read_19_reg_3039_pp0_iter29_reg <= p_read_19_reg_3039_pp0_iter28_reg;
            p_read_19_reg_3039_pp0_iter2_reg <= p_read_19_reg_3039_pp0_iter1_reg;
            p_read_19_reg_3039_pp0_iter30_reg <= p_read_19_reg_3039_pp0_iter29_reg;
            p_read_19_reg_3039_pp0_iter31_reg <= p_read_19_reg_3039_pp0_iter30_reg;
            p_read_19_reg_3039_pp0_iter32_reg <= p_read_19_reg_3039_pp0_iter31_reg;
            p_read_19_reg_3039_pp0_iter33_reg <= p_read_19_reg_3039_pp0_iter32_reg;
            p_read_19_reg_3039_pp0_iter34_reg <= p_read_19_reg_3039_pp0_iter33_reg;
            p_read_19_reg_3039_pp0_iter35_reg <= p_read_19_reg_3039_pp0_iter34_reg;
            p_read_19_reg_3039_pp0_iter36_reg <= p_read_19_reg_3039_pp0_iter35_reg;
            p_read_19_reg_3039_pp0_iter37_reg <= p_read_19_reg_3039_pp0_iter36_reg;
            p_read_19_reg_3039_pp0_iter38_reg <= p_read_19_reg_3039_pp0_iter37_reg;
            p_read_19_reg_3039_pp0_iter39_reg <= p_read_19_reg_3039_pp0_iter38_reg;
            p_read_19_reg_3039_pp0_iter3_reg <= p_read_19_reg_3039_pp0_iter2_reg;
            p_read_19_reg_3039_pp0_iter40_reg <= p_read_19_reg_3039_pp0_iter39_reg;
            p_read_19_reg_3039_pp0_iter41_reg <= p_read_19_reg_3039_pp0_iter40_reg;
            p_read_19_reg_3039_pp0_iter42_reg <= p_read_19_reg_3039_pp0_iter41_reg;
            p_read_19_reg_3039_pp0_iter43_reg <= p_read_19_reg_3039_pp0_iter42_reg;
            p_read_19_reg_3039_pp0_iter44_reg <= p_read_19_reg_3039_pp0_iter43_reg;
            p_read_19_reg_3039_pp0_iter45_reg <= p_read_19_reg_3039_pp0_iter44_reg;
            p_read_19_reg_3039_pp0_iter46_reg <= p_read_19_reg_3039_pp0_iter45_reg;
            p_read_19_reg_3039_pp0_iter47_reg <= p_read_19_reg_3039_pp0_iter46_reg;
            p_read_19_reg_3039_pp0_iter48_reg <= p_read_19_reg_3039_pp0_iter47_reg;
            p_read_19_reg_3039_pp0_iter49_reg <= p_read_19_reg_3039_pp0_iter48_reg;
            p_read_19_reg_3039_pp0_iter4_reg <= p_read_19_reg_3039_pp0_iter3_reg;
            p_read_19_reg_3039_pp0_iter50_reg <= p_read_19_reg_3039_pp0_iter49_reg;
            p_read_19_reg_3039_pp0_iter51_reg <= p_read_19_reg_3039_pp0_iter50_reg;
            p_read_19_reg_3039_pp0_iter52_reg <= p_read_19_reg_3039_pp0_iter51_reg;
            p_read_19_reg_3039_pp0_iter53_reg <= p_read_19_reg_3039_pp0_iter52_reg;
            p_read_19_reg_3039_pp0_iter54_reg <= p_read_19_reg_3039_pp0_iter53_reg;
            p_read_19_reg_3039_pp0_iter55_reg <= p_read_19_reg_3039_pp0_iter54_reg;
            p_read_19_reg_3039_pp0_iter56_reg <= p_read_19_reg_3039_pp0_iter55_reg;
            p_read_19_reg_3039_pp0_iter57_reg <= p_read_19_reg_3039_pp0_iter56_reg;
            p_read_19_reg_3039_pp0_iter58_reg <= p_read_19_reg_3039_pp0_iter57_reg;
            p_read_19_reg_3039_pp0_iter59_reg <= p_read_19_reg_3039_pp0_iter58_reg;
            p_read_19_reg_3039_pp0_iter5_reg <= p_read_19_reg_3039_pp0_iter4_reg;
            p_read_19_reg_3039_pp0_iter60_reg <= p_read_19_reg_3039_pp0_iter59_reg;
            p_read_19_reg_3039_pp0_iter61_reg <= p_read_19_reg_3039_pp0_iter60_reg;
            p_read_19_reg_3039_pp0_iter62_reg <= p_read_19_reg_3039_pp0_iter61_reg;
            p_read_19_reg_3039_pp0_iter63_reg <= p_read_19_reg_3039_pp0_iter62_reg;
            p_read_19_reg_3039_pp0_iter64_reg <= p_read_19_reg_3039_pp0_iter63_reg;
            p_read_19_reg_3039_pp0_iter65_reg <= p_read_19_reg_3039_pp0_iter64_reg;
            p_read_19_reg_3039_pp0_iter66_reg <= p_read_19_reg_3039_pp0_iter65_reg;
            p_read_19_reg_3039_pp0_iter67_reg <= p_read_19_reg_3039_pp0_iter66_reg;
            p_read_19_reg_3039_pp0_iter68_reg <= p_read_19_reg_3039_pp0_iter67_reg;
            p_read_19_reg_3039_pp0_iter69_reg <= p_read_19_reg_3039_pp0_iter68_reg;
            p_read_19_reg_3039_pp0_iter6_reg <= p_read_19_reg_3039_pp0_iter5_reg;
            p_read_19_reg_3039_pp0_iter70_reg <= p_read_19_reg_3039_pp0_iter69_reg;
            p_read_19_reg_3039_pp0_iter71_reg <= p_read_19_reg_3039_pp0_iter70_reg;
            p_read_19_reg_3039_pp0_iter72_reg <= p_read_19_reg_3039_pp0_iter71_reg;
            p_read_19_reg_3039_pp0_iter73_reg <= p_read_19_reg_3039_pp0_iter72_reg;
            p_read_19_reg_3039_pp0_iter74_reg <= p_read_19_reg_3039_pp0_iter73_reg;
            p_read_19_reg_3039_pp0_iter75_reg <= p_read_19_reg_3039_pp0_iter74_reg;
            p_read_19_reg_3039_pp0_iter76_reg <= p_read_19_reg_3039_pp0_iter75_reg;
            p_read_19_reg_3039_pp0_iter7_reg <= p_read_19_reg_3039_pp0_iter6_reg;
            p_read_19_reg_3039_pp0_iter8_reg <= p_read_19_reg_3039_pp0_iter7_reg;
            p_read_19_reg_3039_pp0_iter9_reg <= p_read_19_reg_3039_pp0_iter8_reg;
            p_read_20_reg_3044 <= p_read44_int_reg;
            p_read_20_reg_3044_pp0_iter10_reg <= p_read_20_reg_3044_pp0_iter9_reg;
            p_read_20_reg_3044_pp0_iter11_reg <= p_read_20_reg_3044_pp0_iter10_reg;
            p_read_20_reg_3044_pp0_iter12_reg <= p_read_20_reg_3044_pp0_iter11_reg;
            p_read_20_reg_3044_pp0_iter13_reg <= p_read_20_reg_3044_pp0_iter12_reg;
            p_read_20_reg_3044_pp0_iter14_reg <= p_read_20_reg_3044_pp0_iter13_reg;
            p_read_20_reg_3044_pp0_iter15_reg <= p_read_20_reg_3044_pp0_iter14_reg;
            p_read_20_reg_3044_pp0_iter16_reg <= p_read_20_reg_3044_pp0_iter15_reg;
            p_read_20_reg_3044_pp0_iter17_reg <= p_read_20_reg_3044_pp0_iter16_reg;
            p_read_20_reg_3044_pp0_iter18_reg <= p_read_20_reg_3044_pp0_iter17_reg;
            p_read_20_reg_3044_pp0_iter19_reg <= p_read_20_reg_3044_pp0_iter18_reg;
            p_read_20_reg_3044_pp0_iter1_reg <= p_read_20_reg_3044;
            p_read_20_reg_3044_pp0_iter20_reg <= p_read_20_reg_3044_pp0_iter19_reg;
            p_read_20_reg_3044_pp0_iter21_reg <= p_read_20_reg_3044_pp0_iter20_reg;
            p_read_20_reg_3044_pp0_iter22_reg <= p_read_20_reg_3044_pp0_iter21_reg;
            p_read_20_reg_3044_pp0_iter23_reg <= p_read_20_reg_3044_pp0_iter22_reg;
            p_read_20_reg_3044_pp0_iter24_reg <= p_read_20_reg_3044_pp0_iter23_reg;
            p_read_20_reg_3044_pp0_iter25_reg <= p_read_20_reg_3044_pp0_iter24_reg;
            p_read_20_reg_3044_pp0_iter26_reg <= p_read_20_reg_3044_pp0_iter25_reg;
            p_read_20_reg_3044_pp0_iter27_reg <= p_read_20_reg_3044_pp0_iter26_reg;
            p_read_20_reg_3044_pp0_iter28_reg <= p_read_20_reg_3044_pp0_iter27_reg;
            p_read_20_reg_3044_pp0_iter29_reg <= p_read_20_reg_3044_pp0_iter28_reg;
            p_read_20_reg_3044_pp0_iter2_reg <= p_read_20_reg_3044_pp0_iter1_reg;
            p_read_20_reg_3044_pp0_iter30_reg <= p_read_20_reg_3044_pp0_iter29_reg;
            p_read_20_reg_3044_pp0_iter31_reg <= p_read_20_reg_3044_pp0_iter30_reg;
            p_read_20_reg_3044_pp0_iter32_reg <= p_read_20_reg_3044_pp0_iter31_reg;
            p_read_20_reg_3044_pp0_iter33_reg <= p_read_20_reg_3044_pp0_iter32_reg;
            p_read_20_reg_3044_pp0_iter34_reg <= p_read_20_reg_3044_pp0_iter33_reg;
            p_read_20_reg_3044_pp0_iter35_reg <= p_read_20_reg_3044_pp0_iter34_reg;
            p_read_20_reg_3044_pp0_iter36_reg <= p_read_20_reg_3044_pp0_iter35_reg;
            p_read_20_reg_3044_pp0_iter37_reg <= p_read_20_reg_3044_pp0_iter36_reg;
            p_read_20_reg_3044_pp0_iter38_reg <= p_read_20_reg_3044_pp0_iter37_reg;
            p_read_20_reg_3044_pp0_iter39_reg <= p_read_20_reg_3044_pp0_iter38_reg;
            p_read_20_reg_3044_pp0_iter3_reg <= p_read_20_reg_3044_pp0_iter2_reg;
            p_read_20_reg_3044_pp0_iter40_reg <= p_read_20_reg_3044_pp0_iter39_reg;
            p_read_20_reg_3044_pp0_iter41_reg <= p_read_20_reg_3044_pp0_iter40_reg;
            p_read_20_reg_3044_pp0_iter42_reg <= p_read_20_reg_3044_pp0_iter41_reg;
            p_read_20_reg_3044_pp0_iter43_reg <= p_read_20_reg_3044_pp0_iter42_reg;
            p_read_20_reg_3044_pp0_iter44_reg <= p_read_20_reg_3044_pp0_iter43_reg;
            p_read_20_reg_3044_pp0_iter45_reg <= p_read_20_reg_3044_pp0_iter44_reg;
            p_read_20_reg_3044_pp0_iter46_reg <= p_read_20_reg_3044_pp0_iter45_reg;
            p_read_20_reg_3044_pp0_iter47_reg <= p_read_20_reg_3044_pp0_iter46_reg;
            p_read_20_reg_3044_pp0_iter48_reg <= p_read_20_reg_3044_pp0_iter47_reg;
            p_read_20_reg_3044_pp0_iter49_reg <= p_read_20_reg_3044_pp0_iter48_reg;
            p_read_20_reg_3044_pp0_iter4_reg <= p_read_20_reg_3044_pp0_iter3_reg;
            p_read_20_reg_3044_pp0_iter50_reg <= p_read_20_reg_3044_pp0_iter49_reg;
            p_read_20_reg_3044_pp0_iter51_reg <= p_read_20_reg_3044_pp0_iter50_reg;
            p_read_20_reg_3044_pp0_iter52_reg <= p_read_20_reg_3044_pp0_iter51_reg;
            p_read_20_reg_3044_pp0_iter53_reg <= p_read_20_reg_3044_pp0_iter52_reg;
            p_read_20_reg_3044_pp0_iter54_reg <= p_read_20_reg_3044_pp0_iter53_reg;
            p_read_20_reg_3044_pp0_iter55_reg <= p_read_20_reg_3044_pp0_iter54_reg;
            p_read_20_reg_3044_pp0_iter56_reg <= p_read_20_reg_3044_pp0_iter55_reg;
            p_read_20_reg_3044_pp0_iter57_reg <= p_read_20_reg_3044_pp0_iter56_reg;
            p_read_20_reg_3044_pp0_iter58_reg <= p_read_20_reg_3044_pp0_iter57_reg;
            p_read_20_reg_3044_pp0_iter59_reg <= p_read_20_reg_3044_pp0_iter58_reg;
            p_read_20_reg_3044_pp0_iter5_reg <= p_read_20_reg_3044_pp0_iter4_reg;
            p_read_20_reg_3044_pp0_iter60_reg <= p_read_20_reg_3044_pp0_iter59_reg;
            p_read_20_reg_3044_pp0_iter61_reg <= p_read_20_reg_3044_pp0_iter60_reg;
            p_read_20_reg_3044_pp0_iter62_reg <= p_read_20_reg_3044_pp0_iter61_reg;
            p_read_20_reg_3044_pp0_iter63_reg <= p_read_20_reg_3044_pp0_iter62_reg;
            p_read_20_reg_3044_pp0_iter64_reg <= p_read_20_reg_3044_pp0_iter63_reg;
            p_read_20_reg_3044_pp0_iter65_reg <= p_read_20_reg_3044_pp0_iter64_reg;
            p_read_20_reg_3044_pp0_iter66_reg <= p_read_20_reg_3044_pp0_iter65_reg;
            p_read_20_reg_3044_pp0_iter67_reg <= p_read_20_reg_3044_pp0_iter66_reg;
            p_read_20_reg_3044_pp0_iter68_reg <= p_read_20_reg_3044_pp0_iter67_reg;
            p_read_20_reg_3044_pp0_iter69_reg <= p_read_20_reg_3044_pp0_iter68_reg;
            p_read_20_reg_3044_pp0_iter6_reg <= p_read_20_reg_3044_pp0_iter5_reg;
            p_read_20_reg_3044_pp0_iter70_reg <= p_read_20_reg_3044_pp0_iter69_reg;
            p_read_20_reg_3044_pp0_iter71_reg <= p_read_20_reg_3044_pp0_iter70_reg;
            p_read_20_reg_3044_pp0_iter72_reg <= p_read_20_reg_3044_pp0_iter71_reg;
            p_read_20_reg_3044_pp0_iter73_reg <= p_read_20_reg_3044_pp0_iter72_reg;
            p_read_20_reg_3044_pp0_iter74_reg <= p_read_20_reg_3044_pp0_iter73_reg;
            p_read_20_reg_3044_pp0_iter75_reg <= p_read_20_reg_3044_pp0_iter74_reg;
            p_read_20_reg_3044_pp0_iter76_reg <= p_read_20_reg_3044_pp0_iter75_reg;
            p_read_20_reg_3044_pp0_iter7_reg <= p_read_20_reg_3044_pp0_iter6_reg;
            p_read_20_reg_3044_pp0_iter8_reg <= p_read_20_reg_3044_pp0_iter7_reg;
            p_read_20_reg_3044_pp0_iter9_reg <= p_read_20_reg_3044_pp0_iter8_reg;
            p_read_21_reg_3049 <= p_read43_int_reg;
            p_read_21_reg_3049_pp0_iter10_reg <= p_read_21_reg_3049_pp0_iter9_reg;
            p_read_21_reg_3049_pp0_iter11_reg <= p_read_21_reg_3049_pp0_iter10_reg;
            p_read_21_reg_3049_pp0_iter12_reg <= p_read_21_reg_3049_pp0_iter11_reg;
            p_read_21_reg_3049_pp0_iter13_reg <= p_read_21_reg_3049_pp0_iter12_reg;
            p_read_21_reg_3049_pp0_iter14_reg <= p_read_21_reg_3049_pp0_iter13_reg;
            p_read_21_reg_3049_pp0_iter15_reg <= p_read_21_reg_3049_pp0_iter14_reg;
            p_read_21_reg_3049_pp0_iter16_reg <= p_read_21_reg_3049_pp0_iter15_reg;
            p_read_21_reg_3049_pp0_iter17_reg <= p_read_21_reg_3049_pp0_iter16_reg;
            p_read_21_reg_3049_pp0_iter18_reg <= p_read_21_reg_3049_pp0_iter17_reg;
            p_read_21_reg_3049_pp0_iter19_reg <= p_read_21_reg_3049_pp0_iter18_reg;
            p_read_21_reg_3049_pp0_iter1_reg <= p_read_21_reg_3049;
            p_read_21_reg_3049_pp0_iter20_reg <= p_read_21_reg_3049_pp0_iter19_reg;
            p_read_21_reg_3049_pp0_iter21_reg <= p_read_21_reg_3049_pp0_iter20_reg;
            p_read_21_reg_3049_pp0_iter22_reg <= p_read_21_reg_3049_pp0_iter21_reg;
            p_read_21_reg_3049_pp0_iter23_reg <= p_read_21_reg_3049_pp0_iter22_reg;
            p_read_21_reg_3049_pp0_iter24_reg <= p_read_21_reg_3049_pp0_iter23_reg;
            p_read_21_reg_3049_pp0_iter25_reg <= p_read_21_reg_3049_pp0_iter24_reg;
            p_read_21_reg_3049_pp0_iter26_reg <= p_read_21_reg_3049_pp0_iter25_reg;
            p_read_21_reg_3049_pp0_iter27_reg <= p_read_21_reg_3049_pp0_iter26_reg;
            p_read_21_reg_3049_pp0_iter28_reg <= p_read_21_reg_3049_pp0_iter27_reg;
            p_read_21_reg_3049_pp0_iter29_reg <= p_read_21_reg_3049_pp0_iter28_reg;
            p_read_21_reg_3049_pp0_iter2_reg <= p_read_21_reg_3049_pp0_iter1_reg;
            p_read_21_reg_3049_pp0_iter30_reg <= p_read_21_reg_3049_pp0_iter29_reg;
            p_read_21_reg_3049_pp0_iter31_reg <= p_read_21_reg_3049_pp0_iter30_reg;
            p_read_21_reg_3049_pp0_iter32_reg <= p_read_21_reg_3049_pp0_iter31_reg;
            p_read_21_reg_3049_pp0_iter33_reg <= p_read_21_reg_3049_pp0_iter32_reg;
            p_read_21_reg_3049_pp0_iter34_reg <= p_read_21_reg_3049_pp0_iter33_reg;
            p_read_21_reg_3049_pp0_iter35_reg <= p_read_21_reg_3049_pp0_iter34_reg;
            p_read_21_reg_3049_pp0_iter36_reg <= p_read_21_reg_3049_pp0_iter35_reg;
            p_read_21_reg_3049_pp0_iter37_reg <= p_read_21_reg_3049_pp0_iter36_reg;
            p_read_21_reg_3049_pp0_iter38_reg <= p_read_21_reg_3049_pp0_iter37_reg;
            p_read_21_reg_3049_pp0_iter39_reg <= p_read_21_reg_3049_pp0_iter38_reg;
            p_read_21_reg_3049_pp0_iter3_reg <= p_read_21_reg_3049_pp0_iter2_reg;
            p_read_21_reg_3049_pp0_iter40_reg <= p_read_21_reg_3049_pp0_iter39_reg;
            p_read_21_reg_3049_pp0_iter41_reg <= p_read_21_reg_3049_pp0_iter40_reg;
            p_read_21_reg_3049_pp0_iter42_reg <= p_read_21_reg_3049_pp0_iter41_reg;
            p_read_21_reg_3049_pp0_iter43_reg <= p_read_21_reg_3049_pp0_iter42_reg;
            p_read_21_reg_3049_pp0_iter44_reg <= p_read_21_reg_3049_pp0_iter43_reg;
            p_read_21_reg_3049_pp0_iter45_reg <= p_read_21_reg_3049_pp0_iter44_reg;
            p_read_21_reg_3049_pp0_iter46_reg <= p_read_21_reg_3049_pp0_iter45_reg;
            p_read_21_reg_3049_pp0_iter47_reg <= p_read_21_reg_3049_pp0_iter46_reg;
            p_read_21_reg_3049_pp0_iter48_reg <= p_read_21_reg_3049_pp0_iter47_reg;
            p_read_21_reg_3049_pp0_iter49_reg <= p_read_21_reg_3049_pp0_iter48_reg;
            p_read_21_reg_3049_pp0_iter4_reg <= p_read_21_reg_3049_pp0_iter3_reg;
            p_read_21_reg_3049_pp0_iter50_reg <= p_read_21_reg_3049_pp0_iter49_reg;
            p_read_21_reg_3049_pp0_iter51_reg <= p_read_21_reg_3049_pp0_iter50_reg;
            p_read_21_reg_3049_pp0_iter52_reg <= p_read_21_reg_3049_pp0_iter51_reg;
            p_read_21_reg_3049_pp0_iter53_reg <= p_read_21_reg_3049_pp0_iter52_reg;
            p_read_21_reg_3049_pp0_iter54_reg <= p_read_21_reg_3049_pp0_iter53_reg;
            p_read_21_reg_3049_pp0_iter55_reg <= p_read_21_reg_3049_pp0_iter54_reg;
            p_read_21_reg_3049_pp0_iter56_reg <= p_read_21_reg_3049_pp0_iter55_reg;
            p_read_21_reg_3049_pp0_iter57_reg <= p_read_21_reg_3049_pp0_iter56_reg;
            p_read_21_reg_3049_pp0_iter58_reg <= p_read_21_reg_3049_pp0_iter57_reg;
            p_read_21_reg_3049_pp0_iter59_reg <= p_read_21_reg_3049_pp0_iter58_reg;
            p_read_21_reg_3049_pp0_iter5_reg <= p_read_21_reg_3049_pp0_iter4_reg;
            p_read_21_reg_3049_pp0_iter60_reg <= p_read_21_reg_3049_pp0_iter59_reg;
            p_read_21_reg_3049_pp0_iter61_reg <= p_read_21_reg_3049_pp0_iter60_reg;
            p_read_21_reg_3049_pp0_iter62_reg <= p_read_21_reg_3049_pp0_iter61_reg;
            p_read_21_reg_3049_pp0_iter63_reg <= p_read_21_reg_3049_pp0_iter62_reg;
            p_read_21_reg_3049_pp0_iter64_reg <= p_read_21_reg_3049_pp0_iter63_reg;
            p_read_21_reg_3049_pp0_iter65_reg <= p_read_21_reg_3049_pp0_iter64_reg;
            p_read_21_reg_3049_pp0_iter66_reg <= p_read_21_reg_3049_pp0_iter65_reg;
            p_read_21_reg_3049_pp0_iter67_reg <= p_read_21_reg_3049_pp0_iter66_reg;
            p_read_21_reg_3049_pp0_iter68_reg <= p_read_21_reg_3049_pp0_iter67_reg;
            p_read_21_reg_3049_pp0_iter69_reg <= p_read_21_reg_3049_pp0_iter68_reg;
            p_read_21_reg_3049_pp0_iter6_reg <= p_read_21_reg_3049_pp0_iter5_reg;
            p_read_21_reg_3049_pp0_iter70_reg <= p_read_21_reg_3049_pp0_iter69_reg;
            p_read_21_reg_3049_pp0_iter71_reg <= p_read_21_reg_3049_pp0_iter70_reg;
            p_read_21_reg_3049_pp0_iter72_reg <= p_read_21_reg_3049_pp0_iter71_reg;
            p_read_21_reg_3049_pp0_iter73_reg <= p_read_21_reg_3049_pp0_iter72_reg;
            p_read_21_reg_3049_pp0_iter74_reg <= p_read_21_reg_3049_pp0_iter73_reg;
            p_read_21_reg_3049_pp0_iter75_reg <= p_read_21_reg_3049_pp0_iter74_reg;
            p_read_21_reg_3049_pp0_iter76_reg <= p_read_21_reg_3049_pp0_iter75_reg;
            p_read_21_reg_3049_pp0_iter7_reg <= p_read_21_reg_3049_pp0_iter6_reg;
            p_read_21_reg_3049_pp0_iter8_reg <= p_read_21_reg_3049_pp0_iter7_reg;
            p_read_21_reg_3049_pp0_iter9_reg <= p_read_21_reg_3049_pp0_iter8_reg;
            p_read_22_reg_3054 <= p_read42_int_reg;
            p_read_22_reg_3054_pp0_iter10_reg <= p_read_22_reg_3054_pp0_iter9_reg;
            p_read_22_reg_3054_pp0_iter11_reg <= p_read_22_reg_3054_pp0_iter10_reg;
            p_read_22_reg_3054_pp0_iter12_reg <= p_read_22_reg_3054_pp0_iter11_reg;
            p_read_22_reg_3054_pp0_iter13_reg <= p_read_22_reg_3054_pp0_iter12_reg;
            p_read_22_reg_3054_pp0_iter14_reg <= p_read_22_reg_3054_pp0_iter13_reg;
            p_read_22_reg_3054_pp0_iter15_reg <= p_read_22_reg_3054_pp0_iter14_reg;
            p_read_22_reg_3054_pp0_iter16_reg <= p_read_22_reg_3054_pp0_iter15_reg;
            p_read_22_reg_3054_pp0_iter17_reg <= p_read_22_reg_3054_pp0_iter16_reg;
            p_read_22_reg_3054_pp0_iter18_reg <= p_read_22_reg_3054_pp0_iter17_reg;
            p_read_22_reg_3054_pp0_iter19_reg <= p_read_22_reg_3054_pp0_iter18_reg;
            p_read_22_reg_3054_pp0_iter1_reg <= p_read_22_reg_3054;
            p_read_22_reg_3054_pp0_iter20_reg <= p_read_22_reg_3054_pp0_iter19_reg;
            p_read_22_reg_3054_pp0_iter21_reg <= p_read_22_reg_3054_pp0_iter20_reg;
            p_read_22_reg_3054_pp0_iter22_reg <= p_read_22_reg_3054_pp0_iter21_reg;
            p_read_22_reg_3054_pp0_iter23_reg <= p_read_22_reg_3054_pp0_iter22_reg;
            p_read_22_reg_3054_pp0_iter24_reg <= p_read_22_reg_3054_pp0_iter23_reg;
            p_read_22_reg_3054_pp0_iter25_reg <= p_read_22_reg_3054_pp0_iter24_reg;
            p_read_22_reg_3054_pp0_iter26_reg <= p_read_22_reg_3054_pp0_iter25_reg;
            p_read_22_reg_3054_pp0_iter27_reg <= p_read_22_reg_3054_pp0_iter26_reg;
            p_read_22_reg_3054_pp0_iter28_reg <= p_read_22_reg_3054_pp0_iter27_reg;
            p_read_22_reg_3054_pp0_iter29_reg <= p_read_22_reg_3054_pp0_iter28_reg;
            p_read_22_reg_3054_pp0_iter2_reg <= p_read_22_reg_3054_pp0_iter1_reg;
            p_read_22_reg_3054_pp0_iter30_reg <= p_read_22_reg_3054_pp0_iter29_reg;
            p_read_22_reg_3054_pp0_iter31_reg <= p_read_22_reg_3054_pp0_iter30_reg;
            p_read_22_reg_3054_pp0_iter32_reg <= p_read_22_reg_3054_pp0_iter31_reg;
            p_read_22_reg_3054_pp0_iter33_reg <= p_read_22_reg_3054_pp0_iter32_reg;
            p_read_22_reg_3054_pp0_iter34_reg <= p_read_22_reg_3054_pp0_iter33_reg;
            p_read_22_reg_3054_pp0_iter35_reg <= p_read_22_reg_3054_pp0_iter34_reg;
            p_read_22_reg_3054_pp0_iter36_reg <= p_read_22_reg_3054_pp0_iter35_reg;
            p_read_22_reg_3054_pp0_iter37_reg <= p_read_22_reg_3054_pp0_iter36_reg;
            p_read_22_reg_3054_pp0_iter38_reg <= p_read_22_reg_3054_pp0_iter37_reg;
            p_read_22_reg_3054_pp0_iter39_reg <= p_read_22_reg_3054_pp0_iter38_reg;
            p_read_22_reg_3054_pp0_iter3_reg <= p_read_22_reg_3054_pp0_iter2_reg;
            p_read_22_reg_3054_pp0_iter40_reg <= p_read_22_reg_3054_pp0_iter39_reg;
            p_read_22_reg_3054_pp0_iter41_reg <= p_read_22_reg_3054_pp0_iter40_reg;
            p_read_22_reg_3054_pp0_iter42_reg <= p_read_22_reg_3054_pp0_iter41_reg;
            p_read_22_reg_3054_pp0_iter43_reg <= p_read_22_reg_3054_pp0_iter42_reg;
            p_read_22_reg_3054_pp0_iter44_reg <= p_read_22_reg_3054_pp0_iter43_reg;
            p_read_22_reg_3054_pp0_iter45_reg <= p_read_22_reg_3054_pp0_iter44_reg;
            p_read_22_reg_3054_pp0_iter46_reg <= p_read_22_reg_3054_pp0_iter45_reg;
            p_read_22_reg_3054_pp0_iter47_reg <= p_read_22_reg_3054_pp0_iter46_reg;
            p_read_22_reg_3054_pp0_iter48_reg <= p_read_22_reg_3054_pp0_iter47_reg;
            p_read_22_reg_3054_pp0_iter49_reg <= p_read_22_reg_3054_pp0_iter48_reg;
            p_read_22_reg_3054_pp0_iter4_reg <= p_read_22_reg_3054_pp0_iter3_reg;
            p_read_22_reg_3054_pp0_iter50_reg <= p_read_22_reg_3054_pp0_iter49_reg;
            p_read_22_reg_3054_pp0_iter51_reg <= p_read_22_reg_3054_pp0_iter50_reg;
            p_read_22_reg_3054_pp0_iter52_reg <= p_read_22_reg_3054_pp0_iter51_reg;
            p_read_22_reg_3054_pp0_iter53_reg <= p_read_22_reg_3054_pp0_iter52_reg;
            p_read_22_reg_3054_pp0_iter54_reg <= p_read_22_reg_3054_pp0_iter53_reg;
            p_read_22_reg_3054_pp0_iter55_reg <= p_read_22_reg_3054_pp0_iter54_reg;
            p_read_22_reg_3054_pp0_iter56_reg <= p_read_22_reg_3054_pp0_iter55_reg;
            p_read_22_reg_3054_pp0_iter57_reg <= p_read_22_reg_3054_pp0_iter56_reg;
            p_read_22_reg_3054_pp0_iter58_reg <= p_read_22_reg_3054_pp0_iter57_reg;
            p_read_22_reg_3054_pp0_iter59_reg <= p_read_22_reg_3054_pp0_iter58_reg;
            p_read_22_reg_3054_pp0_iter5_reg <= p_read_22_reg_3054_pp0_iter4_reg;
            p_read_22_reg_3054_pp0_iter60_reg <= p_read_22_reg_3054_pp0_iter59_reg;
            p_read_22_reg_3054_pp0_iter61_reg <= p_read_22_reg_3054_pp0_iter60_reg;
            p_read_22_reg_3054_pp0_iter62_reg <= p_read_22_reg_3054_pp0_iter61_reg;
            p_read_22_reg_3054_pp0_iter63_reg <= p_read_22_reg_3054_pp0_iter62_reg;
            p_read_22_reg_3054_pp0_iter64_reg <= p_read_22_reg_3054_pp0_iter63_reg;
            p_read_22_reg_3054_pp0_iter65_reg <= p_read_22_reg_3054_pp0_iter64_reg;
            p_read_22_reg_3054_pp0_iter66_reg <= p_read_22_reg_3054_pp0_iter65_reg;
            p_read_22_reg_3054_pp0_iter67_reg <= p_read_22_reg_3054_pp0_iter66_reg;
            p_read_22_reg_3054_pp0_iter68_reg <= p_read_22_reg_3054_pp0_iter67_reg;
            p_read_22_reg_3054_pp0_iter69_reg <= p_read_22_reg_3054_pp0_iter68_reg;
            p_read_22_reg_3054_pp0_iter6_reg <= p_read_22_reg_3054_pp0_iter5_reg;
            p_read_22_reg_3054_pp0_iter70_reg <= p_read_22_reg_3054_pp0_iter69_reg;
            p_read_22_reg_3054_pp0_iter71_reg <= p_read_22_reg_3054_pp0_iter70_reg;
            p_read_22_reg_3054_pp0_iter72_reg <= p_read_22_reg_3054_pp0_iter71_reg;
            p_read_22_reg_3054_pp0_iter73_reg <= p_read_22_reg_3054_pp0_iter72_reg;
            p_read_22_reg_3054_pp0_iter74_reg <= p_read_22_reg_3054_pp0_iter73_reg;
            p_read_22_reg_3054_pp0_iter75_reg <= p_read_22_reg_3054_pp0_iter74_reg;
            p_read_22_reg_3054_pp0_iter76_reg <= p_read_22_reg_3054_pp0_iter75_reg;
            p_read_22_reg_3054_pp0_iter7_reg <= p_read_22_reg_3054_pp0_iter6_reg;
            p_read_22_reg_3054_pp0_iter8_reg <= p_read_22_reg_3054_pp0_iter7_reg;
            p_read_22_reg_3054_pp0_iter9_reg <= p_read_22_reg_3054_pp0_iter8_reg;
            p_read_23_reg_3059 <= p_read41_int_reg;
            p_read_23_reg_3059_pp0_iter10_reg <= p_read_23_reg_3059_pp0_iter9_reg;
            p_read_23_reg_3059_pp0_iter11_reg <= p_read_23_reg_3059_pp0_iter10_reg;
            p_read_23_reg_3059_pp0_iter12_reg <= p_read_23_reg_3059_pp0_iter11_reg;
            p_read_23_reg_3059_pp0_iter13_reg <= p_read_23_reg_3059_pp0_iter12_reg;
            p_read_23_reg_3059_pp0_iter14_reg <= p_read_23_reg_3059_pp0_iter13_reg;
            p_read_23_reg_3059_pp0_iter15_reg <= p_read_23_reg_3059_pp0_iter14_reg;
            p_read_23_reg_3059_pp0_iter16_reg <= p_read_23_reg_3059_pp0_iter15_reg;
            p_read_23_reg_3059_pp0_iter17_reg <= p_read_23_reg_3059_pp0_iter16_reg;
            p_read_23_reg_3059_pp0_iter18_reg <= p_read_23_reg_3059_pp0_iter17_reg;
            p_read_23_reg_3059_pp0_iter19_reg <= p_read_23_reg_3059_pp0_iter18_reg;
            p_read_23_reg_3059_pp0_iter1_reg <= p_read_23_reg_3059;
            p_read_23_reg_3059_pp0_iter20_reg <= p_read_23_reg_3059_pp0_iter19_reg;
            p_read_23_reg_3059_pp0_iter21_reg <= p_read_23_reg_3059_pp0_iter20_reg;
            p_read_23_reg_3059_pp0_iter22_reg <= p_read_23_reg_3059_pp0_iter21_reg;
            p_read_23_reg_3059_pp0_iter23_reg <= p_read_23_reg_3059_pp0_iter22_reg;
            p_read_23_reg_3059_pp0_iter24_reg <= p_read_23_reg_3059_pp0_iter23_reg;
            p_read_23_reg_3059_pp0_iter25_reg <= p_read_23_reg_3059_pp0_iter24_reg;
            p_read_23_reg_3059_pp0_iter26_reg <= p_read_23_reg_3059_pp0_iter25_reg;
            p_read_23_reg_3059_pp0_iter27_reg <= p_read_23_reg_3059_pp0_iter26_reg;
            p_read_23_reg_3059_pp0_iter28_reg <= p_read_23_reg_3059_pp0_iter27_reg;
            p_read_23_reg_3059_pp0_iter29_reg <= p_read_23_reg_3059_pp0_iter28_reg;
            p_read_23_reg_3059_pp0_iter2_reg <= p_read_23_reg_3059_pp0_iter1_reg;
            p_read_23_reg_3059_pp0_iter30_reg <= p_read_23_reg_3059_pp0_iter29_reg;
            p_read_23_reg_3059_pp0_iter31_reg <= p_read_23_reg_3059_pp0_iter30_reg;
            p_read_23_reg_3059_pp0_iter32_reg <= p_read_23_reg_3059_pp0_iter31_reg;
            p_read_23_reg_3059_pp0_iter33_reg <= p_read_23_reg_3059_pp0_iter32_reg;
            p_read_23_reg_3059_pp0_iter34_reg <= p_read_23_reg_3059_pp0_iter33_reg;
            p_read_23_reg_3059_pp0_iter35_reg <= p_read_23_reg_3059_pp0_iter34_reg;
            p_read_23_reg_3059_pp0_iter36_reg <= p_read_23_reg_3059_pp0_iter35_reg;
            p_read_23_reg_3059_pp0_iter37_reg <= p_read_23_reg_3059_pp0_iter36_reg;
            p_read_23_reg_3059_pp0_iter38_reg <= p_read_23_reg_3059_pp0_iter37_reg;
            p_read_23_reg_3059_pp0_iter39_reg <= p_read_23_reg_3059_pp0_iter38_reg;
            p_read_23_reg_3059_pp0_iter3_reg <= p_read_23_reg_3059_pp0_iter2_reg;
            p_read_23_reg_3059_pp0_iter40_reg <= p_read_23_reg_3059_pp0_iter39_reg;
            p_read_23_reg_3059_pp0_iter41_reg <= p_read_23_reg_3059_pp0_iter40_reg;
            p_read_23_reg_3059_pp0_iter42_reg <= p_read_23_reg_3059_pp0_iter41_reg;
            p_read_23_reg_3059_pp0_iter43_reg <= p_read_23_reg_3059_pp0_iter42_reg;
            p_read_23_reg_3059_pp0_iter44_reg <= p_read_23_reg_3059_pp0_iter43_reg;
            p_read_23_reg_3059_pp0_iter45_reg <= p_read_23_reg_3059_pp0_iter44_reg;
            p_read_23_reg_3059_pp0_iter46_reg <= p_read_23_reg_3059_pp0_iter45_reg;
            p_read_23_reg_3059_pp0_iter47_reg <= p_read_23_reg_3059_pp0_iter46_reg;
            p_read_23_reg_3059_pp0_iter48_reg <= p_read_23_reg_3059_pp0_iter47_reg;
            p_read_23_reg_3059_pp0_iter49_reg <= p_read_23_reg_3059_pp0_iter48_reg;
            p_read_23_reg_3059_pp0_iter4_reg <= p_read_23_reg_3059_pp0_iter3_reg;
            p_read_23_reg_3059_pp0_iter50_reg <= p_read_23_reg_3059_pp0_iter49_reg;
            p_read_23_reg_3059_pp0_iter51_reg <= p_read_23_reg_3059_pp0_iter50_reg;
            p_read_23_reg_3059_pp0_iter52_reg <= p_read_23_reg_3059_pp0_iter51_reg;
            p_read_23_reg_3059_pp0_iter53_reg <= p_read_23_reg_3059_pp0_iter52_reg;
            p_read_23_reg_3059_pp0_iter54_reg <= p_read_23_reg_3059_pp0_iter53_reg;
            p_read_23_reg_3059_pp0_iter55_reg <= p_read_23_reg_3059_pp0_iter54_reg;
            p_read_23_reg_3059_pp0_iter56_reg <= p_read_23_reg_3059_pp0_iter55_reg;
            p_read_23_reg_3059_pp0_iter57_reg <= p_read_23_reg_3059_pp0_iter56_reg;
            p_read_23_reg_3059_pp0_iter58_reg <= p_read_23_reg_3059_pp0_iter57_reg;
            p_read_23_reg_3059_pp0_iter59_reg <= p_read_23_reg_3059_pp0_iter58_reg;
            p_read_23_reg_3059_pp0_iter5_reg <= p_read_23_reg_3059_pp0_iter4_reg;
            p_read_23_reg_3059_pp0_iter60_reg <= p_read_23_reg_3059_pp0_iter59_reg;
            p_read_23_reg_3059_pp0_iter61_reg <= p_read_23_reg_3059_pp0_iter60_reg;
            p_read_23_reg_3059_pp0_iter62_reg <= p_read_23_reg_3059_pp0_iter61_reg;
            p_read_23_reg_3059_pp0_iter63_reg <= p_read_23_reg_3059_pp0_iter62_reg;
            p_read_23_reg_3059_pp0_iter64_reg <= p_read_23_reg_3059_pp0_iter63_reg;
            p_read_23_reg_3059_pp0_iter65_reg <= p_read_23_reg_3059_pp0_iter64_reg;
            p_read_23_reg_3059_pp0_iter66_reg <= p_read_23_reg_3059_pp0_iter65_reg;
            p_read_23_reg_3059_pp0_iter67_reg <= p_read_23_reg_3059_pp0_iter66_reg;
            p_read_23_reg_3059_pp0_iter68_reg <= p_read_23_reg_3059_pp0_iter67_reg;
            p_read_23_reg_3059_pp0_iter69_reg <= p_read_23_reg_3059_pp0_iter68_reg;
            p_read_23_reg_3059_pp0_iter6_reg <= p_read_23_reg_3059_pp0_iter5_reg;
            p_read_23_reg_3059_pp0_iter70_reg <= p_read_23_reg_3059_pp0_iter69_reg;
            p_read_23_reg_3059_pp0_iter71_reg <= p_read_23_reg_3059_pp0_iter70_reg;
            p_read_23_reg_3059_pp0_iter72_reg <= p_read_23_reg_3059_pp0_iter71_reg;
            p_read_23_reg_3059_pp0_iter73_reg <= p_read_23_reg_3059_pp0_iter72_reg;
            p_read_23_reg_3059_pp0_iter74_reg <= p_read_23_reg_3059_pp0_iter73_reg;
            p_read_23_reg_3059_pp0_iter75_reg <= p_read_23_reg_3059_pp0_iter74_reg;
            p_read_23_reg_3059_pp0_iter76_reg <= p_read_23_reg_3059_pp0_iter75_reg;
            p_read_23_reg_3059_pp0_iter7_reg <= p_read_23_reg_3059_pp0_iter6_reg;
            p_read_23_reg_3059_pp0_iter8_reg <= p_read_23_reg_3059_pp0_iter7_reg;
            p_read_23_reg_3059_pp0_iter9_reg <= p_read_23_reg_3059_pp0_iter8_reg;
            p_read_24_reg_3064 <= p_read40_int_reg;
            p_read_24_reg_3064_pp0_iter10_reg <= p_read_24_reg_3064_pp0_iter9_reg;
            p_read_24_reg_3064_pp0_iter11_reg <= p_read_24_reg_3064_pp0_iter10_reg;
            p_read_24_reg_3064_pp0_iter12_reg <= p_read_24_reg_3064_pp0_iter11_reg;
            p_read_24_reg_3064_pp0_iter13_reg <= p_read_24_reg_3064_pp0_iter12_reg;
            p_read_24_reg_3064_pp0_iter14_reg <= p_read_24_reg_3064_pp0_iter13_reg;
            p_read_24_reg_3064_pp0_iter15_reg <= p_read_24_reg_3064_pp0_iter14_reg;
            p_read_24_reg_3064_pp0_iter16_reg <= p_read_24_reg_3064_pp0_iter15_reg;
            p_read_24_reg_3064_pp0_iter17_reg <= p_read_24_reg_3064_pp0_iter16_reg;
            p_read_24_reg_3064_pp0_iter18_reg <= p_read_24_reg_3064_pp0_iter17_reg;
            p_read_24_reg_3064_pp0_iter19_reg <= p_read_24_reg_3064_pp0_iter18_reg;
            p_read_24_reg_3064_pp0_iter1_reg <= p_read_24_reg_3064;
            p_read_24_reg_3064_pp0_iter20_reg <= p_read_24_reg_3064_pp0_iter19_reg;
            p_read_24_reg_3064_pp0_iter21_reg <= p_read_24_reg_3064_pp0_iter20_reg;
            p_read_24_reg_3064_pp0_iter22_reg <= p_read_24_reg_3064_pp0_iter21_reg;
            p_read_24_reg_3064_pp0_iter23_reg <= p_read_24_reg_3064_pp0_iter22_reg;
            p_read_24_reg_3064_pp0_iter24_reg <= p_read_24_reg_3064_pp0_iter23_reg;
            p_read_24_reg_3064_pp0_iter25_reg <= p_read_24_reg_3064_pp0_iter24_reg;
            p_read_24_reg_3064_pp0_iter26_reg <= p_read_24_reg_3064_pp0_iter25_reg;
            p_read_24_reg_3064_pp0_iter27_reg <= p_read_24_reg_3064_pp0_iter26_reg;
            p_read_24_reg_3064_pp0_iter28_reg <= p_read_24_reg_3064_pp0_iter27_reg;
            p_read_24_reg_3064_pp0_iter29_reg <= p_read_24_reg_3064_pp0_iter28_reg;
            p_read_24_reg_3064_pp0_iter2_reg <= p_read_24_reg_3064_pp0_iter1_reg;
            p_read_24_reg_3064_pp0_iter30_reg <= p_read_24_reg_3064_pp0_iter29_reg;
            p_read_24_reg_3064_pp0_iter31_reg <= p_read_24_reg_3064_pp0_iter30_reg;
            p_read_24_reg_3064_pp0_iter32_reg <= p_read_24_reg_3064_pp0_iter31_reg;
            p_read_24_reg_3064_pp0_iter33_reg <= p_read_24_reg_3064_pp0_iter32_reg;
            p_read_24_reg_3064_pp0_iter34_reg <= p_read_24_reg_3064_pp0_iter33_reg;
            p_read_24_reg_3064_pp0_iter35_reg <= p_read_24_reg_3064_pp0_iter34_reg;
            p_read_24_reg_3064_pp0_iter36_reg <= p_read_24_reg_3064_pp0_iter35_reg;
            p_read_24_reg_3064_pp0_iter37_reg <= p_read_24_reg_3064_pp0_iter36_reg;
            p_read_24_reg_3064_pp0_iter38_reg <= p_read_24_reg_3064_pp0_iter37_reg;
            p_read_24_reg_3064_pp0_iter39_reg <= p_read_24_reg_3064_pp0_iter38_reg;
            p_read_24_reg_3064_pp0_iter3_reg <= p_read_24_reg_3064_pp0_iter2_reg;
            p_read_24_reg_3064_pp0_iter40_reg <= p_read_24_reg_3064_pp0_iter39_reg;
            p_read_24_reg_3064_pp0_iter41_reg <= p_read_24_reg_3064_pp0_iter40_reg;
            p_read_24_reg_3064_pp0_iter42_reg <= p_read_24_reg_3064_pp0_iter41_reg;
            p_read_24_reg_3064_pp0_iter43_reg <= p_read_24_reg_3064_pp0_iter42_reg;
            p_read_24_reg_3064_pp0_iter44_reg <= p_read_24_reg_3064_pp0_iter43_reg;
            p_read_24_reg_3064_pp0_iter45_reg <= p_read_24_reg_3064_pp0_iter44_reg;
            p_read_24_reg_3064_pp0_iter46_reg <= p_read_24_reg_3064_pp0_iter45_reg;
            p_read_24_reg_3064_pp0_iter47_reg <= p_read_24_reg_3064_pp0_iter46_reg;
            p_read_24_reg_3064_pp0_iter48_reg <= p_read_24_reg_3064_pp0_iter47_reg;
            p_read_24_reg_3064_pp0_iter49_reg <= p_read_24_reg_3064_pp0_iter48_reg;
            p_read_24_reg_3064_pp0_iter4_reg <= p_read_24_reg_3064_pp0_iter3_reg;
            p_read_24_reg_3064_pp0_iter50_reg <= p_read_24_reg_3064_pp0_iter49_reg;
            p_read_24_reg_3064_pp0_iter51_reg <= p_read_24_reg_3064_pp0_iter50_reg;
            p_read_24_reg_3064_pp0_iter52_reg <= p_read_24_reg_3064_pp0_iter51_reg;
            p_read_24_reg_3064_pp0_iter53_reg <= p_read_24_reg_3064_pp0_iter52_reg;
            p_read_24_reg_3064_pp0_iter54_reg <= p_read_24_reg_3064_pp0_iter53_reg;
            p_read_24_reg_3064_pp0_iter55_reg <= p_read_24_reg_3064_pp0_iter54_reg;
            p_read_24_reg_3064_pp0_iter56_reg <= p_read_24_reg_3064_pp0_iter55_reg;
            p_read_24_reg_3064_pp0_iter57_reg <= p_read_24_reg_3064_pp0_iter56_reg;
            p_read_24_reg_3064_pp0_iter58_reg <= p_read_24_reg_3064_pp0_iter57_reg;
            p_read_24_reg_3064_pp0_iter59_reg <= p_read_24_reg_3064_pp0_iter58_reg;
            p_read_24_reg_3064_pp0_iter5_reg <= p_read_24_reg_3064_pp0_iter4_reg;
            p_read_24_reg_3064_pp0_iter60_reg <= p_read_24_reg_3064_pp0_iter59_reg;
            p_read_24_reg_3064_pp0_iter61_reg <= p_read_24_reg_3064_pp0_iter60_reg;
            p_read_24_reg_3064_pp0_iter62_reg <= p_read_24_reg_3064_pp0_iter61_reg;
            p_read_24_reg_3064_pp0_iter63_reg <= p_read_24_reg_3064_pp0_iter62_reg;
            p_read_24_reg_3064_pp0_iter64_reg <= p_read_24_reg_3064_pp0_iter63_reg;
            p_read_24_reg_3064_pp0_iter65_reg <= p_read_24_reg_3064_pp0_iter64_reg;
            p_read_24_reg_3064_pp0_iter66_reg <= p_read_24_reg_3064_pp0_iter65_reg;
            p_read_24_reg_3064_pp0_iter67_reg <= p_read_24_reg_3064_pp0_iter66_reg;
            p_read_24_reg_3064_pp0_iter68_reg <= p_read_24_reg_3064_pp0_iter67_reg;
            p_read_24_reg_3064_pp0_iter69_reg <= p_read_24_reg_3064_pp0_iter68_reg;
            p_read_24_reg_3064_pp0_iter6_reg <= p_read_24_reg_3064_pp0_iter5_reg;
            p_read_24_reg_3064_pp0_iter70_reg <= p_read_24_reg_3064_pp0_iter69_reg;
            p_read_24_reg_3064_pp0_iter71_reg <= p_read_24_reg_3064_pp0_iter70_reg;
            p_read_24_reg_3064_pp0_iter72_reg <= p_read_24_reg_3064_pp0_iter71_reg;
            p_read_24_reg_3064_pp0_iter73_reg <= p_read_24_reg_3064_pp0_iter72_reg;
            p_read_24_reg_3064_pp0_iter74_reg <= p_read_24_reg_3064_pp0_iter73_reg;
            p_read_24_reg_3064_pp0_iter75_reg <= p_read_24_reg_3064_pp0_iter74_reg;
            p_read_24_reg_3064_pp0_iter76_reg <= p_read_24_reg_3064_pp0_iter75_reg;
            p_read_24_reg_3064_pp0_iter7_reg <= p_read_24_reg_3064_pp0_iter6_reg;
            p_read_24_reg_3064_pp0_iter8_reg <= p_read_24_reg_3064_pp0_iter7_reg;
            p_read_24_reg_3064_pp0_iter9_reg <= p_read_24_reg_3064_pp0_iter8_reg;
            p_read_25_reg_3069 <= p_read39_int_reg;
            p_read_25_reg_3069_pp0_iter10_reg <= p_read_25_reg_3069_pp0_iter9_reg;
            p_read_25_reg_3069_pp0_iter11_reg <= p_read_25_reg_3069_pp0_iter10_reg;
            p_read_25_reg_3069_pp0_iter12_reg <= p_read_25_reg_3069_pp0_iter11_reg;
            p_read_25_reg_3069_pp0_iter13_reg <= p_read_25_reg_3069_pp0_iter12_reg;
            p_read_25_reg_3069_pp0_iter14_reg <= p_read_25_reg_3069_pp0_iter13_reg;
            p_read_25_reg_3069_pp0_iter15_reg <= p_read_25_reg_3069_pp0_iter14_reg;
            p_read_25_reg_3069_pp0_iter16_reg <= p_read_25_reg_3069_pp0_iter15_reg;
            p_read_25_reg_3069_pp0_iter17_reg <= p_read_25_reg_3069_pp0_iter16_reg;
            p_read_25_reg_3069_pp0_iter18_reg <= p_read_25_reg_3069_pp0_iter17_reg;
            p_read_25_reg_3069_pp0_iter19_reg <= p_read_25_reg_3069_pp0_iter18_reg;
            p_read_25_reg_3069_pp0_iter1_reg <= p_read_25_reg_3069;
            p_read_25_reg_3069_pp0_iter20_reg <= p_read_25_reg_3069_pp0_iter19_reg;
            p_read_25_reg_3069_pp0_iter21_reg <= p_read_25_reg_3069_pp0_iter20_reg;
            p_read_25_reg_3069_pp0_iter22_reg <= p_read_25_reg_3069_pp0_iter21_reg;
            p_read_25_reg_3069_pp0_iter23_reg <= p_read_25_reg_3069_pp0_iter22_reg;
            p_read_25_reg_3069_pp0_iter24_reg <= p_read_25_reg_3069_pp0_iter23_reg;
            p_read_25_reg_3069_pp0_iter25_reg <= p_read_25_reg_3069_pp0_iter24_reg;
            p_read_25_reg_3069_pp0_iter26_reg <= p_read_25_reg_3069_pp0_iter25_reg;
            p_read_25_reg_3069_pp0_iter27_reg <= p_read_25_reg_3069_pp0_iter26_reg;
            p_read_25_reg_3069_pp0_iter28_reg <= p_read_25_reg_3069_pp0_iter27_reg;
            p_read_25_reg_3069_pp0_iter29_reg <= p_read_25_reg_3069_pp0_iter28_reg;
            p_read_25_reg_3069_pp0_iter2_reg <= p_read_25_reg_3069_pp0_iter1_reg;
            p_read_25_reg_3069_pp0_iter30_reg <= p_read_25_reg_3069_pp0_iter29_reg;
            p_read_25_reg_3069_pp0_iter31_reg <= p_read_25_reg_3069_pp0_iter30_reg;
            p_read_25_reg_3069_pp0_iter32_reg <= p_read_25_reg_3069_pp0_iter31_reg;
            p_read_25_reg_3069_pp0_iter33_reg <= p_read_25_reg_3069_pp0_iter32_reg;
            p_read_25_reg_3069_pp0_iter34_reg <= p_read_25_reg_3069_pp0_iter33_reg;
            p_read_25_reg_3069_pp0_iter35_reg <= p_read_25_reg_3069_pp0_iter34_reg;
            p_read_25_reg_3069_pp0_iter36_reg <= p_read_25_reg_3069_pp0_iter35_reg;
            p_read_25_reg_3069_pp0_iter37_reg <= p_read_25_reg_3069_pp0_iter36_reg;
            p_read_25_reg_3069_pp0_iter38_reg <= p_read_25_reg_3069_pp0_iter37_reg;
            p_read_25_reg_3069_pp0_iter39_reg <= p_read_25_reg_3069_pp0_iter38_reg;
            p_read_25_reg_3069_pp0_iter3_reg <= p_read_25_reg_3069_pp0_iter2_reg;
            p_read_25_reg_3069_pp0_iter40_reg <= p_read_25_reg_3069_pp0_iter39_reg;
            p_read_25_reg_3069_pp0_iter41_reg <= p_read_25_reg_3069_pp0_iter40_reg;
            p_read_25_reg_3069_pp0_iter42_reg <= p_read_25_reg_3069_pp0_iter41_reg;
            p_read_25_reg_3069_pp0_iter43_reg <= p_read_25_reg_3069_pp0_iter42_reg;
            p_read_25_reg_3069_pp0_iter44_reg <= p_read_25_reg_3069_pp0_iter43_reg;
            p_read_25_reg_3069_pp0_iter45_reg <= p_read_25_reg_3069_pp0_iter44_reg;
            p_read_25_reg_3069_pp0_iter46_reg <= p_read_25_reg_3069_pp0_iter45_reg;
            p_read_25_reg_3069_pp0_iter47_reg <= p_read_25_reg_3069_pp0_iter46_reg;
            p_read_25_reg_3069_pp0_iter48_reg <= p_read_25_reg_3069_pp0_iter47_reg;
            p_read_25_reg_3069_pp0_iter49_reg <= p_read_25_reg_3069_pp0_iter48_reg;
            p_read_25_reg_3069_pp0_iter4_reg <= p_read_25_reg_3069_pp0_iter3_reg;
            p_read_25_reg_3069_pp0_iter50_reg <= p_read_25_reg_3069_pp0_iter49_reg;
            p_read_25_reg_3069_pp0_iter51_reg <= p_read_25_reg_3069_pp0_iter50_reg;
            p_read_25_reg_3069_pp0_iter52_reg <= p_read_25_reg_3069_pp0_iter51_reg;
            p_read_25_reg_3069_pp0_iter53_reg <= p_read_25_reg_3069_pp0_iter52_reg;
            p_read_25_reg_3069_pp0_iter54_reg <= p_read_25_reg_3069_pp0_iter53_reg;
            p_read_25_reg_3069_pp0_iter55_reg <= p_read_25_reg_3069_pp0_iter54_reg;
            p_read_25_reg_3069_pp0_iter56_reg <= p_read_25_reg_3069_pp0_iter55_reg;
            p_read_25_reg_3069_pp0_iter57_reg <= p_read_25_reg_3069_pp0_iter56_reg;
            p_read_25_reg_3069_pp0_iter58_reg <= p_read_25_reg_3069_pp0_iter57_reg;
            p_read_25_reg_3069_pp0_iter59_reg <= p_read_25_reg_3069_pp0_iter58_reg;
            p_read_25_reg_3069_pp0_iter5_reg <= p_read_25_reg_3069_pp0_iter4_reg;
            p_read_25_reg_3069_pp0_iter60_reg <= p_read_25_reg_3069_pp0_iter59_reg;
            p_read_25_reg_3069_pp0_iter61_reg <= p_read_25_reg_3069_pp0_iter60_reg;
            p_read_25_reg_3069_pp0_iter62_reg <= p_read_25_reg_3069_pp0_iter61_reg;
            p_read_25_reg_3069_pp0_iter63_reg <= p_read_25_reg_3069_pp0_iter62_reg;
            p_read_25_reg_3069_pp0_iter64_reg <= p_read_25_reg_3069_pp0_iter63_reg;
            p_read_25_reg_3069_pp0_iter65_reg <= p_read_25_reg_3069_pp0_iter64_reg;
            p_read_25_reg_3069_pp0_iter66_reg <= p_read_25_reg_3069_pp0_iter65_reg;
            p_read_25_reg_3069_pp0_iter67_reg <= p_read_25_reg_3069_pp0_iter66_reg;
            p_read_25_reg_3069_pp0_iter68_reg <= p_read_25_reg_3069_pp0_iter67_reg;
            p_read_25_reg_3069_pp0_iter69_reg <= p_read_25_reg_3069_pp0_iter68_reg;
            p_read_25_reg_3069_pp0_iter6_reg <= p_read_25_reg_3069_pp0_iter5_reg;
            p_read_25_reg_3069_pp0_iter70_reg <= p_read_25_reg_3069_pp0_iter69_reg;
            p_read_25_reg_3069_pp0_iter71_reg <= p_read_25_reg_3069_pp0_iter70_reg;
            p_read_25_reg_3069_pp0_iter72_reg <= p_read_25_reg_3069_pp0_iter71_reg;
            p_read_25_reg_3069_pp0_iter73_reg <= p_read_25_reg_3069_pp0_iter72_reg;
            p_read_25_reg_3069_pp0_iter74_reg <= p_read_25_reg_3069_pp0_iter73_reg;
            p_read_25_reg_3069_pp0_iter75_reg <= p_read_25_reg_3069_pp0_iter74_reg;
            p_read_25_reg_3069_pp0_iter76_reg <= p_read_25_reg_3069_pp0_iter75_reg;
            p_read_25_reg_3069_pp0_iter7_reg <= p_read_25_reg_3069_pp0_iter6_reg;
            p_read_25_reg_3069_pp0_iter8_reg <= p_read_25_reg_3069_pp0_iter7_reg;
            p_read_25_reg_3069_pp0_iter9_reg <= p_read_25_reg_3069_pp0_iter8_reg;
            p_read_26_reg_3074 <= p_read38_int_reg;
            p_read_26_reg_3074_pp0_iter10_reg <= p_read_26_reg_3074_pp0_iter9_reg;
            p_read_26_reg_3074_pp0_iter11_reg <= p_read_26_reg_3074_pp0_iter10_reg;
            p_read_26_reg_3074_pp0_iter12_reg <= p_read_26_reg_3074_pp0_iter11_reg;
            p_read_26_reg_3074_pp0_iter13_reg <= p_read_26_reg_3074_pp0_iter12_reg;
            p_read_26_reg_3074_pp0_iter14_reg <= p_read_26_reg_3074_pp0_iter13_reg;
            p_read_26_reg_3074_pp0_iter15_reg <= p_read_26_reg_3074_pp0_iter14_reg;
            p_read_26_reg_3074_pp0_iter16_reg <= p_read_26_reg_3074_pp0_iter15_reg;
            p_read_26_reg_3074_pp0_iter17_reg <= p_read_26_reg_3074_pp0_iter16_reg;
            p_read_26_reg_3074_pp0_iter18_reg <= p_read_26_reg_3074_pp0_iter17_reg;
            p_read_26_reg_3074_pp0_iter19_reg <= p_read_26_reg_3074_pp0_iter18_reg;
            p_read_26_reg_3074_pp0_iter1_reg <= p_read_26_reg_3074;
            p_read_26_reg_3074_pp0_iter20_reg <= p_read_26_reg_3074_pp0_iter19_reg;
            p_read_26_reg_3074_pp0_iter21_reg <= p_read_26_reg_3074_pp0_iter20_reg;
            p_read_26_reg_3074_pp0_iter22_reg <= p_read_26_reg_3074_pp0_iter21_reg;
            p_read_26_reg_3074_pp0_iter23_reg <= p_read_26_reg_3074_pp0_iter22_reg;
            p_read_26_reg_3074_pp0_iter24_reg <= p_read_26_reg_3074_pp0_iter23_reg;
            p_read_26_reg_3074_pp0_iter25_reg <= p_read_26_reg_3074_pp0_iter24_reg;
            p_read_26_reg_3074_pp0_iter26_reg <= p_read_26_reg_3074_pp0_iter25_reg;
            p_read_26_reg_3074_pp0_iter27_reg <= p_read_26_reg_3074_pp0_iter26_reg;
            p_read_26_reg_3074_pp0_iter28_reg <= p_read_26_reg_3074_pp0_iter27_reg;
            p_read_26_reg_3074_pp0_iter29_reg <= p_read_26_reg_3074_pp0_iter28_reg;
            p_read_26_reg_3074_pp0_iter2_reg <= p_read_26_reg_3074_pp0_iter1_reg;
            p_read_26_reg_3074_pp0_iter30_reg <= p_read_26_reg_3074_pp0_iter29_reg;
            p_read_26_reg_3074_pp0_iter31_reg <= p_read_26_reg_3074_pp0_iter30_reg;
            p_read_26_reg_3074_pp0_iter32_reg <= p_read_26_reg_3074_pp0_iter31_reg;
            p_read_26_reg_3074_pp0_iter33_reg <= p_read_26_reg_3074_pp0_iter32_reg;
            p_read_26_reg_3074_pp0_iter34_reg <= p_read_26_reg_3074_pp0_iter33_reg;
            p_read_26_reg_3074_pp0_iter35_reg <= p_read_26_reg_3074_pp0_iter34_reg;
            p_read_26_reg_3074_pp0_iter36_reg <= p_read_26_reg_3074_pp0_iter35_reg;
            p_read_26_reg_3074_pp0_iter37_reg <= p_read_26_reg_3074_pp0_iter36_reg;
            p_read_26_reg_3074_pp0_iter38_reg <= p_read_26_reg_3074_pp0_iter37_reg;
            p_read_26_reg_3074_pp0_iter39_reg <= p_read_26_reg_3074_pp0_iter38_reg;
            p_read_26_reg_3074_pp0_iter3_reg <= p_read_26_reg_3074_pp0_iter2_reg;
            p_read_26_reg_3074_pp0_iter40_reg <= p_read_26_reg_3074_pp0_iter39_reg;
            p_read_26_reg_3074_pp0_iter41_reg <= p_read_26_reg_3074_pp0_iter40_reg;
            p_read_26_reg_3074_pp0_iter42_reg <= p_read_26_reg_3074_pp0_iter41_reg;
            p_read_26_reg_3074_pp0_iter43_reg <= p_read_26_reg_3074_pp0_iter42_reg;
            p_read_26_reg_3074_pp0_iter44_reg <= p_read_26_reg_3074_pp0_iter43_reg;
            p_read_26_reg_3074_pp0_iter45_reg <= p_read_26_reg_3074_pp0_iter44_reg;
            p_read_26_reg_3074_pp0_iter46_reg <= p_read_26_reg_3074_pp0_iter45_reg;
            p_read_26_reg_3074_pp0_iter47_reg <= p_read_26_reg_3074_pp0_iter46_reg;
            p_read_26_reg_3074_pp0_iter48_reg <= p_read_26_reg_3074_pp0_iter47_reg;
            p_read_26_reg_3074_pp0_iter49_reg <= p_read_26_reg_3074_pp0_iter48_reg;
            p_read_26_reg_3074_pp0_iter4_reg <= p_read_26_reg_3074_pp0_iter3_reg;
            p_read_26_reg_3074_pp0_iter50_reg <= p_read_26_reg_3074_pp0_iter49_reg;
            p_read_26_reg_3074_pp0_iter51_reg <= p_read_26_reg_3074_pp0_iter50_reg;
            p_read_26_reg_3074_pp0_iter52_reg <= p_read_26_reg_3074_pp0_iter51_reg;
            p_read_26_reg_3074_pp0_iter53_reg <= p_read_26_reg_3074_pp0_iter52_reg;
            p_read_26_reg_3074_pp0_iter54_reg <= p_read_26_reg_3074_pp0_iter53_reg;
            p_read_26_reg_3074_pp0_iter55_reg <= p_read_26_reg_3074_pp0_iter54_reg;
            p_read_26_reg_3074_pp0_iter56_reg <= p_read_26_reg_3074_pp0_iter55_reg;
            p_read_26_reg_3074_pp0_iter57_reg <= p_read_26_reg_3074_pp0_iter56_reg;
            p_read_26_reg_3074_pp0_iter58_reg <= p_read_26_reg_3074_pp0_iter57_reg;
            p_read_26_reg_3074_pp0_iter59_reg <= p_read_26_reg_3074_pp0_iter58_reg;
            p_read_26_reg_3074_pp0_iter5_reg <= p_read_26_reg_3074_pp0_iter4_reg;
            p_read_26_reg_3074_pp0_iter60_reg <= p_read_26_reg_3074_pp0_iter59_reg;
            p_read_26_reg_3074_pp0_iter61_reg <= p_read_26_reg_3074_pp0_iter60_reg;
            p_read_26_reg_3074_pp0_iter62_reg <= p_read_26_reg_3074_pp0_iter61_reg;
            p_read_26_reg_3074_pp0_iter63_reg <= p_read_26_reg_3074_pp0_iter62_reg;
            p_read_26_reg_3074_pp0_iter64_reg <= p_read_26_reg_3074_pp0_iter63_reg;
            p_read_26_reg_3074_pp0_iter65_reg <= p_read_26_reg_3074_pp0_iter64_reg;
            p_read_26_reg_3074_pp0_iter66_reg <= p_read_26_reg_3074_pp0_iter65_reg;
            p_read_26_reg_3074_pp0_iter67_reg <= p_read_26_reg_3074_pp0_iter66_reg;
            p_read_26_reg_3074_pp0_iter68_reg <= p_read_26_reg_3074_pp0_iter67_reg;
            p_read_26_reg_3074_pp0_iter69_reg <= p_read_26_reg_3074_pp0_iter68_reg;
            p_read_26_reg_3074_pp0_iter6_reg <= p_read_26_reg_3074_pp0_iter5_reg;
            p_read_26_reg_3074_pp0_iter70_reg <= p_read_26_reg_3074_pp0_iter69_reg;
            p_read_26_reg_3074_pp0_iter71_reg <= p_read_26_reg_3074_pp0_iter70_reg;
            p_read_26_reg_3074_pp0_iter72_reg <= p_read_26_reg_3074_pp0_iter71_reg;
            p_read_26_reg_3074_pp0_iter73_reg <= p_read_26_reg_3074_pp0_iter72_reg;
            p_read_26_reg_3074_pp0_iter74_reg <= p_read_26_reg_3074_pp0_iter73_reg;
            p_read_26_reg_3074_pp0_iter75_reg <= p_read_26_reg_3074_pp0_iter74_reg;
            p_read_26_reg_3074_pp0_iter76_reg <= p_read_26_reg_3074_pp0_iter75_reg;
            p_read_26_reg_3074_pp0_iter7_reg <= p_read_26_reg_3074_pp0_iter6_reg;
            p_read_26_reg_3074_pp0_iter8_reg <= p_read_26_reg_3074_pp0_iter7_reg;
            p_read_26_reg_3074_pp0_iter9_reg <= p_read_26_reg_3074_pp0_iter8_reg;
            p_read_27_reg_3079 <= p_read37_int_reg;
            p_read_27_reg_3079_pp0_iter10_reg <= p_read_27_reg_3079_pp0_iter9_reg;
            p_read_27_reg_3079_pp0_iter11_reg <= p_read_27_reg_3079_pp0_iter10_reg;
            p_read_27_reg_3079_pp0_iter12_reg <= p_read_27_reg_3079_pp0_iter11_reg;
            p_read_27_reg_3079_pp0_iter13_reg <= p_read_27_reg_3079_pp0_iter12_reg;
            p_read_27_reg_3079_pp0_iter14_reg <= p_read_27_reg_3079_pp0_iter13_reg;
            p_read_27_reg_3079_pp0_iter15_reg <= p_read_27_reg_3079_pp0_iter14_reg;
            p_read_27_reg_3079_pp0_iter16_reg <= p_read_27_reg_3079_pp0_iter15_reg;
            p_read_27_reg_3079_pp0_iter17_reg <= p_read_27_reg_3079_pp0_iter16_reg;
            p_read_27_reg_3079_pp0_iter18_reg <= p_read_27_reg_3079_pp0_iter17_reg;
            p_read_27_reg_3079_pp0_iter19_reg <= p_read_27_reg_3079_pp0_iter18_reg;
            p_read_27_reg_3079_pp0_iter1_reg <= p_read_27_reg_3079;
            p_read_27_reg_3079_pp0_iter20_reg <= p_read_27_reg_3079_pp0_iter19_reg;
            p_read_27_reg_3079_pp0_iter21_reg <= p_read_27_reg_3079_pp0_iter20_reg;
            p_read_27_reg_3079_pp0_iter22_reg <= p_read_27_reg_3079_pp0_iter21_reg;
            p_read_27_reg_3079_pp0_iter23_reg <= p_read_27_reg_3079_pp0_iter22_reg;
            p_read_27_reg_3079_pp0_iter24_reg <= p_read_27_reg_3079_pp0_iter23_reg;
            p_read_27_reg_3079_pp0_iter25_reg <= p_read_27_reg_3079_pp0_iter24_reg;
            p_read_27_reg_3079_pp0_iter26_reg <= p_read_27_reg_3079_pp0_iter25_reg;
            p_read_27_reg_3079_pp0_iter27_reg <= p_read_27_reg_3079_pp0_iter26_reg;
            p_read_27_reg_3079_pp0_iter28_reg <= p_read_27_reg_3079_pp0_iter27_reg;
            p_read_27_reg_3079_pp0_iter29_reg <= p_read_27_reg_3079_pp0_iter28_reg;
            p_read_27_reg_3079_pp0_iter2_reg <= p_read_27_reg_3079_pp0_iter1_reg;
            p_read_27_reg_3079_pp0_iter30_reg <= p_read_27_reg_3079_pp0_iter29_reg;
            p_read_27_reg_3079_pp0_iter31_reg <= p_read_27_reg_3079_pp0_iter30_reg;
            p_read_27_reg_3079_pp0_iter32_reg <= p_read_27_reg_3079_pp0_iter31_reg;
            p_read_27_reg_3079_pp0_iter33_reg <= p_read_27_reg_3079_pp0_iter32_reg;
            p_read_27_reg_3079_pp0_iter34_reg <= p_read_27_reg_3079_pp0_iter33_reg;
            p_read_27_reg_3079_pp0_iter35_reg <= p_read_27_reg_3079_pp0_iter34_reg;
            p_read_27_reg_3079_pp0_iter36_reg <= p_read_27_reg_3079_pp0_iter35_reg;
            p_read_27_reg_3079_pp0_iter37_reg <= p_read_27_reg_3079_pp0_iter36_reg;
            p_read_27_reg_3079_pp0_iter38_reg <= p_read_27_reg_3079_pp0_iter37_reg;
            p_read_27_reg_3079_pp0_iter39_reg <= p_read_27_reg_3079_pp0_iter38_reg;
            p_read_27_reg_3079_pp0_iter3_reg <= p_read_27_reg_3079_pp0_iter2_reg;
            p_read_27_reg_3079_pp0_iter40_reg <= p_read_27_reg_3079_pp0_iter39_reg;
            p_read_27_reg_3079_pp0_iter41_reg <= p_read_27_reg_3079_pp0_iter40_reg;
            p_read_27_reg_3079_pp0_iter42_reg <= p_read_27_reg_3079_pp0_iter41_reg;
            p_read_27_reg_3079_pp0_iter43_reg <= p_read_27_reg_3079_pp0_iter42_reg;
            p_read_27_reg_3079_pp0_iter44_reg <= p_read_27_reg_3079_pp0_iter43_reg;
            p_read_27_reg_3079_pp0_iter45_reg <= p_read_27_reg_3079_pp0_iter44_reg;
            p_read_27_reg_3079_pp0_iter46_reg <= p_read_27_reg_3079_pp0_iter45_reg;
            p_read_27_reg_3079_pp0_iter47_reg <= p_read_27_reg_3079_pp0_iter46_reg;
            p_read_27_reg_3079_pp0_iter48_reg <= p_read_27_reg_3079_pp0_iter47_reg;
            p_read_27_reg_3079_pp0_iter49_reg <= p_read_27_reg_3079_pp0_iter48_reg;
            p_read_27_reg_3079_pp0_iter4_reg <= p_read_27_reg_3079_pp0_iter3_reg;
            p_read_27_reg_3079_pp0_iter50_reg <= p_read_27_reg_3079_pp0_iter49_reg;
            p_read_27_reg_3079_pp0_iter51_reg <= p_read_27_reg_3079_pp0_iter50_reg;
            p_read_27_reg_3079_pp0_iter52_reg <= p_read_27_reg_3079_pp0_iter51_reg;
            p_read_27_reg_3079_pp0_iter53_reg <= p_read_27_reg_3079_pp0_iter52_reg;
            p_read_27_reg_3079_pp0_iter54_reg <= p_read_27_reg_3079_pp0_iter53_reg;
            p_read_27_reg_3079_pp0_iter55_reg <= p_read_27_reg_3079_pp0_iter54_reg;
            p_read_27_reg_3079_pp0_iter56_reg <= p_read_27_reg_3079_pp0_iter55_reg;
            p_read_27_reg_3079_pp0_iter57_reg <= p_read_27_reg_3079_pp0_iter56_reg;
            p_read_27_reg_3079_pp0_iter58_reg <= p_read_27_reg_3079_pp0_iter57_reg;
            p_read_27_reg_3079_pp0_iter59_reg <= p_read_27_reg_3079_pp0_iter58_reg;
            p_read_27_reg_3079_pp0_iter5_reg <= p_read_27_reg_3079_pp0_iter4_reg;
            p_read_27_reg_3079_pp0_iter60_reg <= p_read_27_reg_3079_pp0_iter59_reg;
            p_read_27_reg_3079_pp0_iter61_reg <= p_read_27_reg_3079_pp0_iter60_reg;
            p_read_27_reg_3079_pp0_iter62_reg <= p_read_27_reg_3079_pp0_iter61_reg;
            p_read_27_reg_3079_pp0_iter63_reg <= p_read_27_reg_3079_pp0_iter62_reg;
            p_read_27_reg_3079_pp0_iter64_reg <= p_read_27_reg_3079_pp0_iter63_reg;
            p_read_27_reg_3079_pp0_iter65_reg <= p_read_27_reg_3079_pp0_iter64_reg;
            p_read_27_reg_3079_pp0_iter66_reg <= p_read_27_reg_3079_pp0_iter65_reg;
            p_read_27_reg_3079_pp0_iter67_reg <= p_read_27_reg_3079_pp0_iter66_reg;
            p_read_27_reg_3079_pp0_iter68_reg <= p_read_27_reg_3079_pp0_iter67_reg;
            p_read_27_reg_3079_pp0_iter69_reg <= p_read_27_reg_3079_pp0_iter68_reg;
            p_read_27_reg_3079_pp0_iter6_reg <= p_read_27_reg_3079_pp0_iter5_reg;
            p_read_27_reg_3079_pp0_iter70_reg <= p_read_27_reg_3079_pp0_iter69_reg;
            p_read_27_reg_3079_pp0_iter71_reg <= p_read_27_reg_3079_pp0_iter70_reg;
            p_read_27_reg_3079_pp0_iter72_reg <= p_read_27_reg_3079_pp0_iter71_reg;
            p_read_27_reg_3079_pp0_iter73_reg <= p_read_27_reg_3079_pp0_iter72_reg;
            p_read_27_reg_3079_pp0_iter74_reg <= p_read_27_reg_3079_pp0_iter73_reg;
            p_read_27_reg_3079_pp0_iter75_reg <= p_read_27_reg_3079_pp0_iter74_reg;
            p_read_27_reg_3079_pp0_iter76_reg <= p_read_27_reg_3079_pp0_iter75_reg;
            p_read_27_reg_3079_pp0_iter7_reg <= p_read_27_reg_3079_pp0_iter6_reg;
            p_read_27_reg_3079_pp0_iter8_reg <= p_read_27_reg_3079_pp0_iter7_reg;
            p_read_27_reg_3079_pp0_iter9_reg <= p_read_27_reg_3079_pp0_iter8_reg;
            p_read_28_reg_3084 <= p_read36_int_reg;
            p_read_28_reg_3084_pp0_iter10_reg <= p_read_28_reg_3084_pp0_iter9_reg;
            p_read_28_reg_3084_pp0_iter11_reg <= p_read_28_reg_3084_pp0_iter10_reg;
            p_read_28_reg_3084_pp0_iter12_reg <= p_read_28_reg_3084_pp0_iter11_reg;
            p_read_28_reg_3084_pp0_iter13_reg <= p_read_28_reg_3084_pp0_iter12_reg;
            p_read_28_reg_3084_pp0_iter14_reg <= p_read_28_reg_3084_pp0_iter13_reg;
            p_read_28_reg_3084_pp0_iter15_reg <= p_read_28_reg_3084_pp0_iter14_reg;
            p_read_28_reg_3084_pp0_iter16_reg <= p_read_28_reg_3084_pp0_iter15_reg;
            p_read_28_reg_3084_pp0_iter17_reg <= p_read_28_reg_3084_pp0_iter16_reg;
            p_read_28_reg_3084_pp0_iter18_reg <= p_read_28_reg_3084_pp0_iter17_reg;
            p_read_28_reg_3084_pp0_iter19_reg <= p_read_28_reg_3084_pp0_iter18_reg;
            p_read_28_reg_3084_pp0_iter1_reg <= p_read_28_reg_3084;
            p_read_28_reg_3084_pp0_iter20_reg <= p_read_28_reg_3084_pp0_iter19_reg;
            p_read_28_reg_3084_pp0_iter21_reg <= p_read_28_reg_3084_pp0_iter20_reg;
            p_read_28_reg_3084_pp0_iter22_reg <= p_read_28_reg_3084_pp0_iter21_reg;
            p_read_28_reg_3084_pp0_iter23_reg <= p_read_28_reg_3084_pp0_iter22_reg;
            p_read_28_reg_3084_pp0_iter24_reg <= p_read_28_reg_3084_pp0_iter23_reg;
            p_read_28_reg_3084_pp0_iter25_reg <= p_read_28_reg_3084_pp0_iter24_reg;
            p_read_28_reg_3084_pp0_iter26_reg <= p_read_28_reg_3084_pp0_iter25_reg;
            p_read_28_reg_3084_pp0_iter27_reg <= p_read_28_reg_3084_pp0_iter26_reg;
            p_read_28_reg_3084_pp0_iter28_reg <= p_read_28_reg_3084_pp0_iter27_reg;
            p_read_28_reg_3084_pp0_iter29_reg <= p_read_28_reg_3084_pp0_iter28_reg;
            p_read_28_reg_3084_pp0_iter2_reg <= p_read_28_reg_3084_pp0_iter1_reg;
            p_read_28_reg_3084_pp0_iter30_reg <= p_read_28_reg_3084_pp0_iter29_reg;
            p_read_28_reg_3084_pp0_iter31_reg <= p_read_28_reg_3084_pp0_iter30_reg;
            p_read_28_reg_3084_pp0_iter32_reg <= p_read_28_reg_3084_pp0_iter31_reg;
            p_read_28_reg_3084_pp0_iter33_reg <= p_read_28_reg_3084_pp0_iter32_reg;
            p_read_28_reg_3084_pp0_iter34_reg <= p_read_28_reg_3084_pp0_iter33_reg;
            p_read_28_reg_3084_pp0_iter35_reg <= p_read_28_reg_3084_pp0_iter34_reg;
            p_read_28_reg_3084_pp0_iter36_reg <= p_read_28_reg_3084_pp0_iter35_reg;
            p_read_28_reg_3084_pp0_iter37_reg <= p_read_28_reg_3084_pp0_iter36_reg;
            p_read_28_reg_3084_pp0_iter38_reg <= p_read_28_reg_3084_pp0_iter37_reg;
            p_read_28_reg_3084_pp0_iter39_reg <= p_read_28_reg_3084_pp0_iter38_reg;
            p_read_28_reg_3084_pp0_iter3_reg <= p_read_28_reg_3084_pp0_iter2_reg;
            p_read_28_reg_3084_pp0_iter40_reg <= p_read_28_reg_3084_pp0_iter39_reg;
            p_read_28_reg_3084_pp0_iter41_reg <= p_read_28_reg_3084_pp0_iter40_reg;
            p_read_28_reg_3084_pp0_iter42_reg <= p_read_28_reg_3084_pp0_iter41_reg;
            p_read_28_reg_3084_pp0_iter43_reg <= p_read_28_reg_3084_pp0_iter42_reg;
            p_read_28_reg_3084_pp0_iter44_reg <= p_read_28_reg_3084_pp0_iter43_reg;
            p_read_28_reg_3084_pp0_iter45_reg <= p_read_28_reg_3084_pp0_iter44_reg;
            p_read_28_reg_3084_pp0_iter46_reg <= p_read_28_reg_3084_pp0_iter45_reg;
            p_read_28_reg_3084_pp0_iter47_reg <= p_read_28_reg_3084_pp0_iter46_reg;
            p_read_28_reg_3084_pp0_iter48_reg <= p_read_28_reg_3084_pp0_iter47_reg;
            p_read_28_reg_3084_pp0_iter49_reg <= p_read_28_reg_3084_pp0_iter48_reg;
            p_read_28_reg_3084_pp0_iter4_reg <= p_read_28_reg_3084_pp0_iter3_reg;
            p_read_28_reg_3084_pp0_iter50_reg <= p_read_28_reg_3084_pp0_iter49_reg;
            p_read_28_reg_3084_pp0_iter51_reg <= p_read_28_reg_3084_pp0_iter50_reg;
            p_read_28_reg_3084_pp0_iter52_reg <= p_read_28_reg_3084_pp0_iter51_reg;
            p_read_28_reg_3084_pp0_iter53_reg <= p_read_28_reg_3084_pp0_iter52_reg;
            p_read_28_reg_3084_pp0_iter54_reg <= p_read_28_reg_3084_pp0_iter53_reg;
            p_read_28_reg_3084_pp0_iter55_reg <= p_read_28_reg_3084_pp0_iter54_reg;
            p_read_28_reg_3084_pp0_iter56_reg <= p_read_28_reg_3084_pp0_iter55_reg;
            p_read_28_reg_3084_pp0_iter57_reg <= p_read_28_reg_3084_pp0_iter56_reg;
            p_read_28_reg_3084_pp0_iter58_reg <= p_read_28_reg_3084_pp0_iter57_reg;
            p_read_28_reg_3084_pp0_iter59_reg <= p_read_28_reg_3084_pp0_iter58_reg;
            p_read_28_reg_3084_pp0_iter5_reg <= p_read_28_reg_3084_pp0_iter4_reg;
            p_read_28_reg_3084_pp0_iter60_reg <= p_read_28_reg_3084_pp0_iter59_reg;
            p_read_28_reg_3084_pp0_iter61_reg <= p_read_28_reg_3084_pp0_iter60_reg;
            p_read_28_reg_3084_pp0_iter62_reg <= p_read_28_reg_3084_pp0_iter61_reg;
            p_read_28_reg_3084_pp0_iter63_reg <= p_read_28_reg_3084_pp0_iter62_reg;
            p_read_28_reg_3084_pp0_iter64_reg <= p_read_28_reg_3084_pp0_iter63_reg;
            p_read_28_reg_3084_pp0_iter65_reg <= p_read_28_reg_3084_pp0_iter64_reg;
            p_read_28_reg_3084_pp0_iter66_reg <= p_read_28_reg_3084_pp0_iter65_reg;
            p_read_28_reg_3084_pp0_iter67_reg <= p_read_28_reg_3084_pp0_iter66_reg;
            p_read_28_reg_3084_pp0_iter68_reg <= p_read_28_reg_3084_pp0_iter67_reg;
            p_read_28_reg_3084_pp0_iter69_reg <= p_read_28_reg_3084_pp0_iter68_reg;
            p_read_28_reg_3084_pp0_iter6_reg <= p_read_28_reg_3084_pp0_iter5_reg;
            p_read_28_reg_3084_pp0_iter70_reg <= p_read_28_reg_3084_pp0_iter69_reg;
            p_read_28_reg_3084_pp0_iter71_reg <= p_read_28_reg_3084_pp0_iter70_reg;
            p_read_28_reg_3084_pp0_iter72_reg <= p_read_28_reg_3084_pp0_iter71_reg;
            p_read_28_reg_3084_pp0_iter73_reg <= p_read_28_reg_3084_pp0_iter72_reg;
            p_read_28_reg_3084_pp0_iter74_reg <= p_read_28_reg_3084_pp0_iter73_reg;
            p_read_28_reg_3084_pp0_iter75_reg <= p_read_28_reg_3084_pp0_iter74_reg;
            p_read_28_reg_3084_pp0_iter76_reg <= p_read_28_reg_3084_pp0_iter75_reg;
            p_read_28_reg_3084_pp0_iter7_reg <= p_read_28_reg_3084_pp0_iter6_reg;
            p_read_28_reg_3084_pp0_iter8_reg <= p_read_28_reg_3084_pp0_iter7_reg;
            p_read_28_reg_3084_pp0_iter9_reg <= p_read_28_reg_3084_pp0_iter8_reg;
            p_read_29_reg_3089 <= p_read35_int_reg;
            p_read_29_reg_3089_pp0_iter10_reg <= p_read_29_reg_3089_pp0_iter9_reg;
            p_read_29_reg_3089_pp0_iter11_reg <= p_read_29_reg_3089_pp0_iter10_reg;
            p_read_29_reg_3089_pp0_iter12_reg <= p_read_29_reg_3089_pp0_iter11_reg;
            p_read_29_reg_3089_pp0_iter13_reg <= p_read_29_reg_3089_pp0_iter12_reg;
            p_read_29_reg_3089_pp0_iter14_reg <= p_read_29_reg_3089_pp0_iter13_reg;
            p_read_29_reg_3089_pp0_iter15_reg <= p_read_29_reg_3089_pp0_iter14_reg;
            p_read_29_reg_3089_pp0_iter16_reg <= p_read_29_reg_3089_pp0_iter15_reg;
            p_read_29_reg_3089_pp0_iter17_reg <= p_read_29_reg_3089_pp0_iter16_reg;
            p_read_29_reg_3089_pp0_iter18_reg <= p_read_29_reg_3089_pp0_iter17_reg;
            p_read_29_reg_3089_pp0_iter19_reg <= p_read_29_reg_3089_pp0_iter18_reg;
            p_read_29_reg_3089_pp0_iter1_reg <= p_read_29_reg_3089;
            p_read_29_reg_3089_pp0_iter20_reg <= p_read_29_reg_3089_pp0_iter19_reg;
            p_read_29_reg_3089_pp0_iter21_reg <= p_read_29_reg_3089_pp0_iter20_reg;
            p_read_29_reg_3089_pp0_iter22_reg <= p_read_29_reg_3089_pp0_iter21_reg;
            p_read_29_reg_3089_pp0_iter23_reg <= p_read_29_reg_3089_pp0_iter22_reg;
            p_read_29_reg_3089_pp0_iter24_reg <= p_read_29_reg_3089_pp0_iter23_reg;
            p_read_29_reg_3089_pp0_iter25_reg <= p_read_29_reg_3089_pp0_iter24_reg;
            p_read_29_reg_3089_pp0_iter26_reg <= p_read_29_reg_3089_pp0_iter25_reg;
            p_read_29_reg_3089_pp0_iter27_reg <= p_read_29_reg_3089_pp0_iter26_reg;
            p_read_29_reg_3089_pp0_iter28_reg <= p_read_29_reg_3089_pp0_iter27_reg;
            p_read_29_reg_3089_pp0_iter29_reg <= p_read_29_reg_3089_pp0_iter28_reg;
            p_read_29_reg_3089_pp0_iter2_reg <= p_read_29_reg_3089_pp0_iter1_reg;
            p_read_29_reg_3089_pp0_iter30_reg <= p_read_29_reg_3089_pp0_iter29_reg;
            p_read_29_reg_3089_pp0_iter31_reg <= p_read_29_reg_3089_pp0_iter30_reg;
            p_read_29_reg_3089_pp0_iter32_reg <= p_read_29_reg_3089_pp0_iter31_reg;
            p_read_29_reg_3089_pp0_iter33_reg <= p_read_29_reg_3089_pp0_iter32_reg;
            p_read_29_reg_3089_pp0_iter34_reg <= p_read_29_reg_3089_pp0_iter33_reg;
            p_read_29_reg_3089_pp0_iter35_reg <= p_read_29_reg_3089_pp0_iter34_reg;
            p_read_29_reg_3089_pp0_iter36_reg <= p_read_29_reg_3089_pp0_iter35_reg;
            p_read_29_reg_3089_pp0_iter37_reg <= p_read_29_reg_3089_pp0_iter36_reg;
            p_read_29_reg_3089_pp0_iter38_reg <= p_read_29_reg_3089_pp0_iter37_reg;
            p_read_29_reg_3089_pp0_iter39_reg <= p_read_29_reg_3089_pp0_iter38_reg;
            p_read_29_reg_3089_pp0_iter3_reg <= p_read_29_reg_3089_pp0_iter2_reg;
            p_read_29_reg_3089_pp0_iter40_reg <= p_read_29_reg_3089_pp0_iter39_reg;
            p_read_29_reg_3089_pp0_iter41_reg <= p_read_29_reg_3089_pp0_iter40_reg;
            p_read_29_reg_3089_pp0_iter42_reg <= p_read_29_reg_3089_pp0_iter41_reg;
            p_read_29_reg_3089_pp0_iter43_reg <= p_read_29_reg_3089_pp0_iter42_reg;
            p_read_29_reg_3089_pp0_iter44_reg <= p_read_29_reg_3089_pp0_iter43_reg;
            p_read_29_reg_3089_pp0_iter45_reg <= p_read_29_reg_3089_pp0_iter44_reg;
            p_read_29_reg_3089_pp0_iter46_reg <= p_read_29_reg_3089_pp0_iter45_reg;
            p_read_29_reg_3089_pp0_iter47_reg <= p_read_29_reg_3089_pp0_iter46_reg;
            p_read_29_reg_3089_pp0_iter48_reg <= p_read_29_reg_3089_pp0_iter47_reg;
            p_read_29_reg_3089_pp0_iter49_reg <= p_read_29_reg_3089_pp0_iter48_reg;
            p_read_29_reg_3089_pp0_iter4_reg <= p_read_29_reg_3089_pp0_iter3_reg;
            p_read_29_reg_3089_pp0_iter50_reg <= p_read_29_reg_3089_pp0_iter49_reg;
            p_read_29_reg_3089_pp0_iter51_reg <= p_read_29_reg_3089_pp0_iter50_reg;
            p_read_29_reg_3089_pp0_iter52_reg <= p_read_29_reg_3089_pp0_iter51_reg;
            p_read_29_reg_3089_pp0_iter53_reg <= p_read_29_reg_3089_pp0_iter52_reg;
            p_read_29_reg_3089_pp0_iter54_reg <= p_read_29_reg_3089_pp0_iter53_reg;
            p_read_29_reg_3089_pp0_iter55_reg <= p_read_29_reg_3089_pp0_iter54_reg;
            p_read_29_reg_3089_pp0_iter56_reg <= p_read_29_reg_3089_pp0_iter55_reg;
            p_read_29_reg_3089_pp0_iter57_reg <= p_read_29_reg_3089_pp0_iter56_reg;
            p_read_29_reg_3089_pp0_iter58_reg <= p_read_29_reg_3089_pp0_iter57_reg;
            p_read_29_reg_3089_pp0_iter59_reg <= p_read_29_reg_3089_pp0_iter58_reg;
            p_read_29_reg_3089_pp0_iter5_reg <= p_read_29_reg_3089_pp0_iter4_reg;
            p_read_29_reg_3089_pp0_iter60_reg <= p_read_29_reg_3089_pp0_iter59_reg;
            p_read_29_reg_3089_pp0_iter61_reg <= p_read_29_reg_3089_pp0_iter60_reg;
            p_read_29_reg_3089_pp0_iter62_reg <= p_read_29_reg_3089_pp0_iter61_reg;
            p_read_29_reg_3089_pp0_iter63_reg <= p_read_29_reg_3089_pp0_iter62_reg;
            p_read_29_reg_3089_pp0_iter64_reg <= p_read_29_reg_3089_pp0_iter63_reg;
            p_read_29_reg_3089_pp0_iter65_reg <= p_read_29_reg_3089_pp0_iter64_reg;
            p_read_29_reg_3089_pp0_iter66_reg <= p_read_29_reg_3089_pp0_iter65_reg;
            p_read_29_reg_3089_pp0_iter67_reg <= p_read_29_reg_3089_pp0_iter66_reg;
            p_read_29_reg_3089_pp0_iter68_reg <= p_read_29_reg_3089_pp0_iter67_reg;
            p_read_29_reg_3089_pp0_iter69_reg <= p_read_29_reg_3089_pp0_iter68_reg;
            p_read_29_reg_3089_pp0_iter6_reg <= p_read_29_reg_3089_pp0_iter5_reg;
            p_read_29_reg_3089_pp0_iter70_reg <= p_read_29_reg_3089_pp0_iter69_reg;
            p_read_29_reg_3089_pp0_iter71_reg <= p_read_29_reg_3089_pp0_iter70_reg;
            p_read_29_reg_3089_pp0_iter72_reg <= p_read_29_reg_3089_pp0_iter71_reg;
            p_read_29_reg_3089_pp0_iter73_reg <= p_read_29_reg_3089_pp0_iter72_reg;
            p_read_29_reg_3089_pp0_iter74_reg <= p_read_29_reg_3089_pp0_iter73_reg;
            p_read_29_reg_3089_pp0_iter75_reg <= p_read_29_reg_3089_pp0_iter74_reg;
            p_read_29_reg_3089_pp0_iter76_reg <= p_read_29_reg_3089_pp0_iter75_reg;
            p_read_29_reg_3089_pp0_iter7_reg <= p_read_29_reg_3089_pp0_iter6_reg;
            p_read_29_reg_3089_pp0_iter8_reg <= p_read_29_reg_3089_pp0_iter7_reg;
            p_read_29_reg_3089_pp0_iter9_reg <= p_read_29_reg_3089_pp0_iter8_reg;
            p_read_30_reg_3094 <= p_read34_int_reg;
            p_read_30_reg_3094_pp0_iter10_reg <= p_read_30_reg_3094_pp0_iter9_reg;
            p_read_30_reg_3094_pp0_iter11_reg <= p_read_30_reg_3094_pp0_iter10_reg;
            p_read_30_reg_3094_pp0_iter12_reg <= p_read_30_reg_3094_pp0_iter11_reg;
            p_read_30_reg_3094_pp0_iter13_reg <= p_read_30_reg_3094_pp0_iter12_reg;
            p_read_30_reg_3094_pp0_iter14_reg <= p_read_30_reg_3094_pp0_iter13_reg;
            p_read_30_reg_3094_pp0_iter15_reg <= p_read_30_reg_3094_pp0_iter14_reg;
            p_read_30_reg_3094_pp0_iter16_reg <= p_read_30_reg_3094_pp0_iter15_reg;
            p_read_30_reg_3094_pp0_iter17_reg <= p_read_30_reg_3094_pp0_iter16_reg;
            p_read_30_reg_3094_pp0_iter18_reg <= p_read_30_reg_3094_pp0_iter17_reg;
            p_read_30_reg_3094_pp0_iter19_reg <= p_read_30_reg_3094_pp0_iter18_reg;
            p_read_30_reg_3094_pp0_iter1_reg <= p_read_30_reg_3094;
            p_read_30_reg_3094_pp0_iter20_reg <= p_read_30_reg_3094_pp0_iter19_reg;
            p_read_30_reg_3094_pp0_iter21_reg <= p_read_30_reg_3094_pp0_iter20_reg;
            p_read_30_reg_3094_pp0_iter22_reg <= p_read_30_reg_3094_pp0_iter21_reg;
            p_read_30_reg_3094_pp0_iter23_reg <= p_read_30_reg_3094_pp0_iter22_reg;
            p_read_30_reg_3094_pp0_iter24_reg <= p_read_30_reg_3094_pp0_iter23_reg;
            p_read_30_reg_3094_pp0_iter25_reg <= p_read_30_reg_3094_pp0_iter24_reg;
            p_read_30_reg_3094_pp0_iter26_reg <= p_read_30_reg_3094_pp0_iter25_reg;
            p_read_30_reg_3094_pp0_iter27_reg <= p_read_30_reg_3094_pp0_iter26_reg;
            p_read_30_reg_3094_pp0_iter28_reg <= p_read_30_reg_3094_pp0_iter27_reg;
            p_read_30_reg_3094_pp0_iter29_reg <= p_read_30_reg_3094_pp0_iter28_reg;
            p_read_30_reg_3094_pp0_iter2_reg <= p_read_30_reg_3094_pp0_iter1_reg;
            p_read_30_reg_3094_pp0_iter30_reg <= p_read_30_reg_3094_pp0_iter29_reg;
            p_read_30_reg_3094_pp0_iter31_reg <= p_read_30_reg_3094_pp0_iter30_reg;
            p_read_30_reg_3094_pp0_iter32_reg <= p_read_30_reg_3094_pp0_iter31_reg;
            p_read_30_reg_3094_pp0_iter33_reg <= p_read_30_reg_3094_pp0_iter32_reg;
            p_read_30_reg_3094_pp0_iter34_reg <= p_read_30_reg_3094_pp0_iter33_reg;
            p_read_30_reg_3094_pp0_iter35_reg <= p_read_30_reg_3094_pp0_iter34_reg;
            p_read_30_reg_3094_pp0_iter36_reg <= p_read_30_reg_3094_pp0_iter35_reg;
            p_read_30_reg_3094_pp0_iter37_reg <= p_read_30_reg_3094_pp0_iter36_reg;
            p_read_30_reg_3094_pp0_iter38_reg <= p_read_30_reg_3094_pp0_iter37_reg;
            p_read_30_reg_3094_pp0_iter39_reg <= p_read_30_reg_3094_pp0_iter38_reg;
            p_read_30_reg_3094_pp0_iter3_reg <= p_read_30_reg_3094_pp0_iter2_reg;
            p_read_30_reg_3094_pp0_iter40_reg <= p_read_30_reg_3094_pp0_iter39_reg;
            p_read_30_reg_3094_pp0_iter41_reg <= p_read_30_reg_3094_pp0_iter40_reg;
            p_read_30_reg_3094_pp0_iter42_reg <= p_read_30_reg_3094_pp0_iter41_reg;
            p_read_30_reg_3094_pp0_iter43_reg <= p_read_30_reg_3094_pp0_iter42_reg;
            p_read_30_reg_3094_pp0_iter44_reg <= p_read_30_reg_3094_pp0_iter43_reg;
            p_read_30_reg_3094_pp0_iter45_reg <= p_read_30_reg_3094_pp0_iter44_reg;
            p_read_30_reg_3094_pp0_iter46_reg <= p_read_30_reg_3094_pp0_iter45_reg;
            p_read_30_reg_3094_pp0_iter47_reg <= p_read_30_reg_3094_pp0_iter46_reg;
            p_read_30_reg_3094_pp0_iter48_reg <= p_read_30_reg_3094_pp0_iter47_reg;
            p_read_30_reg_3094_pp0_iter49_reg <= p_read_30_reg_3094_pp0_iter48_reg;
            p_read_30_reg_3094_pp0_iter4_reg <= p_read_30_reg_3094_pp0_iter3_reg;
            p_read_30_reg_3094_pp0_iter50_reg <= p_read_30_reg_3094_pp0_iter49_reg;
            p_read_30_reg_3094_pp0_iter51_reg <= p_read_30_reg_3094_pp0_iter50_reg;
            p_read_30_reg_3094_pp0_iter52_reg <= p_read_30_reg_3094_pp0_iter51_reg;
            p_read_30_reg_3094_pp0_iter53_reg <= p_read_30_reg_3094_pp0_iter52_reg;
            p_read_30_reg_3094_pp0_iter54_reg <= p_read_30_reg_3094_pp0_iter53_reg;
            p_read_30_reg_3094_pp0_iter55_reg <= p_read_30_reg_3094_pp0_iter54_reg;
            p_read_30_reg_3094_pp0_iter56_reg <= p_read_30_reg_3094_pp0_iter55_reg;
            p_read_30_reg_3094_pp0_iter57_reg <= p_read_30_reg_3094_pp0_iter56_reg;
            p_read_30_reg_3094_pp0_iter58_reg <= p_read_30_reg_3094_pp0_iter57_reg;
            p_read_30_reg_3094_pp0_iter59_reg <= p_read_30_reg_3094_pp0_iter58_reg;
            p_read_30_reg_3094_pp0_iter5_reg <= p_read_30_reg_3094_pp0_iter4_reg;
            p_read_30_reg_3094_pp0_iter60_reg <= p_read_30_reg_3094_pp0_iter59_reg;
            p_read_30_reg_3094_pp0_iter61_reg <= p_read_30_reg_3094_pp0_iter60_reg;
            p_read_30_reg_3094_pp0_iter62_reg <= p_read_30_reg_3094_pp0_iter61_reg;
            p_read_30_reg_3094_pp0_iter63_reg <= p_read_30_reg_3094_pp0_iter62_reg;
            p_read_30_reg_3094_pp0_iter64_reg <= p_read_30_reg_3094_pp0_iter63_reg;
            p_read_30_reg_3094_pp0_iter65_reg <= p_read_30_reg_3094_pp0_iter64_reg;
            p_read_30_reg_3094_pp0_iter66_reg <= p_read_30_reg_3094_pp0_iter65_reg;
            p_read_30_reg_3094_pp0_iter67_reg <= p_read_30_reg_3094_pp0_iter66_reg;
            p_read_30_reg_3094_pp0_iter68_reg <= p_read_30_reg_3094_pp0_iter67_reg;
            p_read_30_reg_3094_pp0_iter69_reg <= p_read_30_reg_3094_pp0_iter68_reg;
            p_read_30_reg_3094_pp0_iter6_reg <= p_read_30_reg_3094_pp0_iter5_reg;
            p_read_30_reg_3094_pp0_iter70_reg <= p_read_30_reg_3094_pp0_iter69_reg;
            p_read_30_reg_3094_pp0_iter71_reg <= p_read_30_reg_3094_pp0_iter70_reg;
            p_read_30_reg_3094_pp0_iter72_reg <= p_read_30_reg_3094_pp0_iter71_reg;
            p_read_30_reg_3094_pp0_iter73_reg <= p_read_30_reg_3094_pp0_iter72_reg;
            p_read_30_reg_3094_pp0_iter74_reg <= p_read_30_reg_3094_pp0_iter73_reg;
            p_read_30_reg_3094_pp0_iter75_reg <= p_read_30_reg_3094_pp0_iter74_reg;
            p_read_30_reg_3094_pp0_iter76_reg <= p_read_30_reg_3094_pp0_iter75_reg;
            p_read_30_reg_3094_pp0_iter7_reg <= p_read_30_reg_3094_pp0_iter6_reg;
            p_read_30_reg_3094_pp0_iter8_reg <= p_read_30_reg_3094_pp0_iter7_reg;
            p_read_30_reg_3094_pp0_iter9_reg <= p_read_30_reg_3094_pp0_iter8_reg;
            p_read_31_reg_3099 <= p_read33_int_reg;
            p_read_31_reg_3099_pp0_iter10_reg <= p_read_31_reg_3099_pp0_iter9_reg;
            p_read_31_reg_3099_pp0_iter11_reg <= p_read_31_reg_3099_pp0_iter10_reg;
            p_read_31_reg_3099_pp0_iter12_reg <= p_read_31_reg_3099_pp0_iter11_reg;
            p_read_31_reg_3099_pp0_iter13_reg <= p_read_31_reg_3099_pp0_iter12_reg;
            p_read_31_reg_3099_pp0_iter14_reg <= p_read_31_reg_3099_pp0_iter13_reg;
            p_read_31_reg_3099_pp0_iter15_reg <= p_read_31_reg_3099_pp0_iter14_reg;
            p_read_31_reg_3099_pp0_iter16_reg <= p_read_31_reg_3099_pp0_iter15_reg;
            p_read_31_reg_3099_pp0_iter17_reg <= p_read_31_reg_3099_pp0_iter16_reg;
            p_read_31_reg_3099_pp0_iter18_reg <= p_read_31_reg_3099_pp0_iter17_reg;
            p_read_31_reg_3099_pp0_iter19_reg <= p_read_31_reg_3099_pp0_iter18_reg;
            p_read_31_reg_3099_pp0_iter1_reg <= p_read_31_reg_3099;
            p_read_31_reg_3099_pp0_iter20_reg <= p_read_31_reg_3099_pp0_iter19_reg;
            p_read_31_reg_3099_pp0_iter21_reg <= p_read_31_reg_3099_pp0_iter20_reg;
            p_read_31_reg_3099_pp0_iter22_reg <= p_read_31_reg_3099_pp0_iter21_reg;
            p_read_31_reg_3099_pp0_iter23_reg <= p_read_31_reg_3099_pp0_iter22_reg;
            p_read_31_reg_3099_pp0_iter24_reg <= p_read_31_reg_3099_pp0_iter23_reg;
            p_read_31_reg_3099_pp0_iter25_reg <= p_read_31_reg_3099_pp0_iter24_reg;
            p_read_31_reg_3099_pp0_iter26_reg <= p_read_31_reg_3099_pp0_iter25_reg;
            p_read_31_reg_3099_pp0_iter27_reg <= p_read_31_reg_3099_pp0_iter26_reg;
            p_read_31_reg_3099_pp0_iter28_reg <= p_read_31_reg_3099_pp0_iter27_reg;
            p_read_31_reg_3099_pp0_iter29_reg <= p_read_31_reg_3099_pp0_iter28_reg;
            p_read_31_reg_3099_pp0_iter2_reg <= p_read_31_reg_3099_pp0_iter1_reg;
            p_read_31_reg_3099_pp0_iter30_reg <= p_read_31_reg_3099_pp0_iter29_reg;
            p_read_31_reg_3099_pp0_iter31_reg <= p_read_31_reg_3099_pp0_iter30_reg;
            p_read_31_reg_3099_pp0_iter32_reg <= p_read_31_reg_3099_pp0_iter31_reg;
            p_read_31_reg_3099_pp0_iter33_reg <= p_read_31_reg_3099_pp0_iter32_reg;
            p_read_31_reg_3099_pp0_iter34_reg <= p_read_31_reg_3099_pp0_iter33_reg;
            p_read_31_reg_3099_pp0_iter35_reg <= p_read_31_reg_3099_pp0_iter34_reg;
            p_read_31_reg_3099_pp0_iter36_reg <= p_read_31_reg_3099_pp0_iter35_reg;
            p_read_31_reg_3099_pp0_iter37_reg <= p_read_31_reg_3099_pp0_iter36_reg;
            p_read_31_reg_3099_pp0_iter38_reg <= p_read_31_reg_3099_pp0_iter37_reg;
            p_read_31_reg_3099_pp0_iter39_reg <= p_read_31_reg_3099_pp0_iter38_reg;
            p_read_31_reg_3099_pp0_iter3_reg <= p_read_31_reg_3099_pp0_iter2_reg;
            p_read_31_reg_3099_pp0_iter40_reg <= p_read_31_reg_3099_pp0_iter39_reg;
            p_read_31_reg_3099_pp0_iter41_reg <= p_read_31_reg_3099_pp0_iter40_reg;
            p_read_31_reg_3099_pp0_iter42_reg <= p_read_31_reg_3099_pp0_iter41_reg;
            p_read_31_reg_3099_pp0_iter43_reg <= p_read_31_reg_3099_pp0_iter42_reg;
            p_read_31_reg_3099_pp0_iter44_reg <= p_read_31_reg_3099_pp0_iter43_reg;
            p_read_31_reg_3099_pp0_iter45_reg <= p_read_31_reg_3099_pp0_iter44_reg;
            p_read_31_reg_3099_pp0_iter46_reg <= p_read_31_reg_3099_pp0_iter45_reg;
            p_read_31_reg_3099_pp0_iter47_reg <= p_read_31_reg_3099_pp0_iter46_reg;
            p_read_31_reg_3099_pp0_iter48_reg <= p_read_31_reg_3099_pp0_iter47_reg;
            p_read_31_reg_3099_pp0_iter49_reg <= p_read_31_reg_3099_pp0_iter48_reg;
            p_read_31_reg_3099_pp0_iter4_reg <= p_read_31_reg_3099_pp0_iter3_reg;
            p_read_31_reg_3099_pp0_iter50_reg <= p_read_31_reg_3099_pp0_iter49_reg;
            p_read_31_reg_3099_pp0_iter51_reg <= p_read_31_reg_3099_pp0_iter50_reg;
            p_read_31_reg_3099_pp0_iter52_reg <= p_read_31_reg_3099_pp0_iter51_reg;
            p_read_31_reg_3099_pp0_iter53_reg <= p_read_31_reg_3099_pp0_iter52_reg;
            p_read_31_reg_3099_pp0_iter54_reg <= p_read_31_reg_3099_pp0_iter53_reg;
            p_read_31_reg_3099_pp0_iter55_reg <= p_read_31_reg_3099_pp0_iter54_reg;
            p_read_31_reg_3099_pp0_iter56_reg <= p_read_31_reg_3099_pp0_iter55_reg;
            p_read_31_reg_3099_pp0_iter57_reg <= p_read_31_reg_3099_pp0_iter56_reg;
            p_read_31_reg_3099_pp0_iter58_reg <= p_read_31_reg_3099_pp0_iter57_reg;
            p_read_31_reg_3099_pp0_iter59_reg <= p_read_31_reg_3099_pp0_iter58_reg;
            p_read_31_reg_3099_pp0_iter5_reg <= p_read_31_reg_3099_pp0_iter4_reg;
            p_read_31_reg_3099_pp0_iter60_reg <= p_read_31_reg_3099_pp0_iter59_reg;
            p_read_31_reg_3099_pp0_iter61_reg <= p_read_31_reg_3099_pp0_iter60_reg;
            p_read_31_reg_3099_pp0_iter62_reg <= p_read_31_reg_3099_pp0_iter61_reg;
            p_read_31_reg_3099_pp0_iter63_reg <= p_read_31_reg_3099_pp0_iter62_reg;
            p_read_31_reg_3099_pp0_iter64_reg <= p_read_31_reg_3099_pp0_iter63_reg;
            p_read_31_reg_3099_pp0_iter65_reg <= p_read_31_reg_3099_pp0_iter64_reg;
            p_read_31_reg_3099_pp0_iter66_reg <= p_read_31_reg_3099_pp0_iter65_reg;
            p_read_31_reg_3099_pp0_iter67_reg <= p_read_31_reg_3099_pp0_iter66_reg;
            p_read_31_reg_3099_pp0_iter68_reg <= p_read_31_reg_3099_pp0_iter67_reg;
            p_read_31_reg_3099_pp0_iter69_reg <= p_read_31_reg_3099_pp0_iter68_reg;
            p_read_31_reg_3099_pp0_iter6_reg <= p_read_31_reg_3099_pp0_iter5_reg;
            p_read_31_reg_3099_pp0_iter70_reg <= p_read_31_reg_3099_pp0_iter69_reg;
            p_read_31_reg_3099_pp0_iter71_reg <= p_read_31_reg_3099_pp0_iter70_reg;
            p_read_31_reg_3099_pp0_iter72_reg <= p_read_31_reg_3099_pp0_iter71_reg;
            p_read_31_reg_3099_pp0_iter73_reg <= p_read_31_reg_3099_pp0_iter72_reg;
            p_read_31_reg_3099_pp0_iter74_reg <= p_read_31_reg_3099_pp0_iter73_reg;
            p_read_31_reg_3099_pp0_iter75_reg <= p_read_31_reg_3099_pp0_iter74_reg;
            p_read_31_reg_3099_pp0_iter76_reg <= p_read_31_reg_3099_pp0_iter75_reg;
            p_read_31_reg_3099_pp0_iter7_reg <= p_read_31_reg_3099_pp0_iter6_reg;
            p_read_31_reg_3099_pp0_iter8_reg <= p_read_31_reg_3099_pp0_iter7_reg;
            p_read_31_reg_3099_pp0_iter9_reg <= p_read_31_reg_3099_pp0_iter8_reg;
            p_read_32_reg_3104 <= p_read32_int_reg;
            p_read_32_reg_3104_pp0_iter10_reg <= p_read_32_reg_3104_pp0_iter9_reg;
            p_read_32_reg_3104_pp0_iter11_reg <= p_read_32_reg_3104_pp0_iter10_reg;
            p_read_32_reg_3104_pp0_iter12_reg <= p_read_32_reg_3104_pp0_iter11_reg;
            p_read_32_reg_3104_pp0_iter13_reg <= p_read_32_reg_3104_pp0_iter12_reg;
            p_read_32_reg_3104_pp0_iter14_reg <= p_read_32_reg_3104_pp0_iter13_reg;
            p_read_32_reg_3104_pp0_iter15_reg <= p_read_32_reg_3104_pp0_iter14_reg;
            p_read_32_reg_3104_pp0_iter16_reg <= p_read_32_reg_3104_pp0_iter15_reg;
            p_read_32_reg_3104_pp0_iter17_reg <= p_read_32_reg_3104_pp0_iter16_reg;
            p_read_32_reg_3104_pp0_iter18_reg <= p_read_32_reg_3104_pp0_iter17_reg;
            p_read_32_reg_3104_pp0_iter19_reg <= p_read_32_reg_3104_pp0_iter18_reg;
            p_read_32_reg_3104_pp0_iter1_reg <= p_read_32_reg_3104;
            p_read_32_reg_3104_pp0_iter20_reg <= p_read_32_reg_3104_pp0_iter19_reg;
            p_read_32_reg_3104_pp0_iter21_reg <= p_read_32_reg_3104_pp0_iter20_reg;
            p_read_32_reg_3104_pp0_iter22_reg <= p_read_32_reg_3104_pp0_iter21_reg;
            p_read_32_reg_3104_pp0_iter23_reg <= p_read_32_reg_3104_pp0_iter22_reg;
            p_read_32_reg_3104_pp0_iter24_reg <= p_read_32_reg_3104_pp0_iter23_reg;
            p_read_32_reg_3104_pp0_iter25_reg <= p_read_32_reg_3104_pp0_iter24_reg;
            p_read_32_reg_3104_pp0_iter26_reg <= p_read_32_reg_3104_pp0_iter25_reg;
            p_read_32_reg_3104_pp0_iter27_reg <= p_read_32_reg_3104_pp0_iter26_reg;
            p_read_32_reg_3104_pp0_iter28_reg <= p_read_32_reg_3104_pp0_iter27_reg;
            p_read_32_reg_3104_pp0_iter29_reg <= p_read_32_reg_3104_pp0_iter28_reg;
            p_read_32_reg_3104_pp0_iter2_reg <= p_read_32_reg_3104_pp0_iter1_reg;
            p_read_32_reg_3104_pp0_iter30_reg <= p_read_32_reg_3104_pp0_iter29_reg;
            p_read_32_reg_3104_pp0_iter31_reg <= p_read_32_reg_3104_pp0_iter30_reg;
            p_read_32_reg_3104_pp0_iter32_reg <= p_read_32_reg_3104_pp0_iter31_reg;
            p_read_32_reg_3104_pp0_iter33_reg <= p_read_32_reg_3104_pp0_iter32_reg;
            p_read_32_reg_3104_pp0_iter34_reg <= p_read_32_reg_3104_pp0_iter33_reg;
            p_read_32_reg_3104_pp0_iter35_reg <= p_read_32_reg_3104_pp0_iter34_reg;
            p_read_32_reg_3104_pp0_iter36_reg <= p_read_32_reg_3104_pp0_iter35_reg;
            p_read_32_reg_3104_pp0_iter37_reg <= p_read_32_reg_3104_pp0_iter36_reg;
            p_read_32_reg_3104_pp0_iter38_reg <= p_read_32_reg_3104_pp0_iter37_reg;
            p_read_32_reg_3104_pp0_iter39_reg <= p_read_32_reg_3104_pp0_iter38_reg;
            p_read_32_reg_3104_pp0_iter3_reg <= p_read_32_reg_3104_pp0_iter2_reg;
            p_read_32_reg_3104_pp0_iter40_reg <= p_read_32_reg_3104_pp0_iter39_reg;
            p_read_32_reg_3104_pp0_iter41_reg <= p_read_32_reg_3104_pp0_iter40_reg;
            p_read_32_reg_3104_pp0_iter42_reg <= p_read_32_reg_3104_pp0_iter41_reg;
            p_read_32_reg_3104_pp0_iter43_reg <= p_read_32_reg_3104_pp0_iter42_reg;
            p_read_32_reg_3104_pp0_iter44_reg <= p_read_32_reg_3104_pp0_iter43_reg;
            p_read_32_reg_3104_pp0_iter45_reg <= p_read_32_reg_3104_pp0_iter44_reg;
            p_read_32_reg_3104_pp0_iter46_reg <= p_read_32_reg_3104_pp0_iter45_reg;
            p_read_32_reg_3104_pp0_iter47_reg <= p_read_32_reg_3104_pp0_iter46_reg;
            p_read_32_reg_3104_pp0_iter48_reg <= p_read_32_reg_3104_pp0_iter47_reg;
            p_read_32_reg_3104_pp0_iter49_reg <= p_read_32_reg_3104_pp0_iter48_reg;
            p_read_32_reg_3104_pp0_iter4_reg <= p_read_32_reg_3104_pp0_iter3_reg;
            p_read_32_reg_3104_pp0_iter50_reg <= p_read_32_reg_3104_pp0_iter49_reg;
            p_read_32_reg_3104_pp0_iter51_reg <= p_read_32_reg_3104_pp0_iter50_reg;
            p_read_32_reg_3104_pp0_iter52_reg <= p_read_32_reg_3104_pp0_iter51_reg;
            p_read_32_reg_3104_pp0_iter53_reg <= p_read_32_reg_3104_pp0_iter52_reg;
            p_read_32_reg_3104_pp0_iter54_reg <= p_read_32_reg_3104_pp0_iter53_reg;
            p_read_32_reg_3104_pp0_iter55_reg <= p_read_32_reg_3104_pp0_iter54_reg;
            p_read_32_reg_3104_pp0_iter56_reg <= p_read_32_reg_3104_pp0_iter55_reg;
            p_read_32_reg_3104_pp0_iter57_reg <= p_read_32_reg_3104_pp0_iter56_reg;
            p_read_32_reg_3104_pp0_iter58_reg <= p_read_32_reg_3104_pp0_iter57_reg;
            p_read_32_reg_3104_pp0_iter59_reg <= p_read_32_reg_3104_pp0_iter58_reg;
            p_read_32_reg_3104_pp0_iter5_reg <= p_read_32_reg_3104_pp0_iter4_reg;
            p_read_32_reg_3104_pp0_iter60_reg <= p_read_32_reg_3104_pp0_iter59_reg;
            p_read_32_reg_3104_pp0_iter61_reg <= p_read_32_reg_3104_pp0_iter60_reg;
            p_read_32_reg_3104_pp0_iter62_reg <= p_read_32_reg_3104_pp0_iter61_reg;
            p_read_32_reg_3104_pp0_iter63_reg <= p_read_32_reg_3104_pp0_iter62_reg;
            p_read_32_reg_3104_pp0_iter64_reg <= p_read_32_reg_3104_pp0_iter63_reg;
            p_read_32_reg_3104_pp0_iter65_reg <= p_read_32_reg_3104_pp0_iter64_reg;
            p_read_32_reg_3104_pp0_iter66_reg <= p_read_32_reg_3104_pp0_iter65_reg;
            p_read_32_reg_3104_pp0_iter67_reg <= p_read_32_reg_3104_pp0_iter66_reg;
            p_read_32_reg_3104_pp0_iter68_reg <= p_read_32_reg_3104_pp0_iter67_reg;
            p_read_32_reg_3104_pp0_iter69_reg <= p_read_32_reg_3104_pp0_iter68_reg;
            p_read_32_reg_3104_pp0_iter6_reg <= p_read_32_reg_3104_pp0_iter5_reg;
            p_read_32_reg_3104_pp0_iter70_reg <= p_read_32_reg_3104_pp0_iter69_reg;
            p_read_32_reg_3104_pp0_iter71_reg <= p_read_32_reg_3104_pp0_iter70_reg;
            p_read_32_reg_3104_pp0_iter72_reg <= p_read_32_reg_3104_pp0_iter71_reg;
            p_read_32_reg_3104_pp0_iter73_reg <= p_read_32_reg_3104_pp0_iter72_reg;
            p_read_32_reg_3104_pp0_iter74_reg <= p_read_32_reg_3104_pp0_iter73_reg;
            p_read_32_reg_3104_pp0_iter75_reg <= p_read_32_reg_3104_pp0_iter74_reg;
            p_read_32_reg_3104_pp0_iter76_reg <= p_read_32_reg_3104_pp0_iter75_reg;
            p_read_32_reg_3104_pp0_iter7_reg <= p_read_32_reg_3104_pp0_iter6_reg;
            p_read_32_reg_3104_pp0_iter8_reg <= p_read_32_reg_3104_pp0_iter7_reg;
            p_read_32_reg_3104_pp0_iter9_reg <= p_read_32_reg_3104_pp0_iter8_reg;
            p_read_33_reg_3109 <= p_read31_int_reg;
            p_read_33_reg_3109_pp0_iter10_reg <= p_read_33_reg_3109_pp0_iter9_reg;
            p_read_33_reg_3109_pp0_iter11_reg <= p_read_33_reg_3109_pp0_iter10_reg;
            p_read_33_reg_3109_pp0_iter12_reg <= p_read_33_reg_3109_pp0_iter11_reg;
            p_read_33_reg_3109_pp0_iter13_reg <= p_read_33_reg_3109_pp0_iter12_reg;
            p_read_33_reg_3109_pp0_iter14_reg <= p_read_33_reg_3109_pp0_iter13_reg;
            p_read_33_reg_3109_pp0_iter15_reg <= p_read_33_reg_3109_pp0_iter14_reg;
            p_read_33_reg_3109_pp0_iter16_reg <= p_read_33_reg_3109_pp0_iter15_reg;
            p_read_33_reg_3109_pp0_iter17_reg <= p_read_33_reg_3109_pp0_iter16_reg;
            p_read_33_reg_3109_pp0_iter18_reg <= p_read_33_reg_3109_pp0_iter17_reg;
            p_read_33_reg_3109_pp0_iter19_reg <= p_read_33_reg_3109_pp0_iter18_reg;
            p_read_33_reg_3109_pp0_iter1_reg <= p_read_33_reg_3109;
            p_read_33_reg_3109_pp0_iter20_reg <= p_read_33_reg_3109_pp0_iter19_reg;
            p_read_33_reg_3109_pp0_iter21_reg <= p_read_33_reg_3109_pp0_iter20_reg;
            p_read_33_reg_3109_pp0_iter22_reg <= p_read_33_reg_3109_pp0_iter21_reg;
            p_read_33_reg_3109_pp0_iter23_reg <= p_read_33_reg_3109_pp0_iter22_reg;
            p_read_33_reg_3109_pp0_iter24_reg <= p_read_33_reg_3109_pp0_iter23_reg;
            p_read_33_reg_3109_pp0_iter25_reg <= p_read_33_reg_3109_pp0_iter24_reg;
            p_read_33_reg_3109_pp0_iter26_reg <= p_read_33_reg_3109_pp0_iter25_reg;
            p_read_33_reg_3109_pp0_iter27_reg <= p_read_33_reg_3109_pp0_iter26_reg;
            p_read_33_reg_3109_pp0_iter28_reg <= p_read_33_reg_3109_pp0_iter27_reg;
            p_read_33_reg_3109_pp0_iter29_reg <= p_read_33_reg_3109_pp0_iter28_reg;
            p_read_33_reg_3109_pp0_iter2_reg <= p_read_33_reg_3109_pp0_iter1_reg;
            p_read_33_reg_3109_pp0_iter30_reg <= p_read_33_reg_3109_pp0_iter29_reg;
            p_read_33_reg_3109_pp0_iter31_reg <= p_read_33_reg_3109_pp0_iter30_reg;
            p_read_33_reg_3109_pp0_iter32_reg <= p_read_33_reg_3109_pp0_iter31_reg;
            p_read_33_reg_3109_pp0_iter33_reg <= p_read_33_reg_3109_pp0_iter32_reg;
            p_read_33_reg_3109_pp0_iter34_reg <= p_read_33_reg_3109_pp0_iter33_reg;
            p_read_33_reg_3109_pp0_iter35_reg <= p_read_33_reg_3109_pp0_iter34_reg;
            p_read_33_reg_3109_pp0_iter36_reg <= p_read_33_reg_3109_pp0_iter35_reg;
            p_read_33_reg_3109_pp0_iter37_reg <= p_read_33_reg_3109_pp0_iter36_reg;
            p_read_33_reg_3109_pp0_iter38_reg <= p_read_33_reg_3109_pp0_iter37_reg;
            p_read_33_reg_3109_pp0_iter39_reg <= p_read_33_reg_3109_pp0_iter38_reg;
            p_read_33_reg_3109_pp0_iter3_reg <= p_read_33_reg_3109_pp0_iter2_reg;
            p_read_33_reg_3109_pp0_iter40_reg <= p_read_33_reg_3109_pp0_iter39_reg;
            p_read_33_reg_3109_pp0_iter41_reg <= p_read_33_reg_3109_pp0_iter40_reg;
            p_read_33_reg_3109_pp0_iter42_reg <= p_read_33_reg_3109_pp0_iter41_reg;
            p_read_33_reg_3109_pp0_iter43_reg <= p_read_33_reg_3109_pp0_iter42_reg;
            p_read_33_reg_3109_pp0_iter44_reg <= p_read_33_reg_3109_pp0_iter43_reg;
            p_read_33_reg_3109_pp0_iter45_reg <= p_read_33_reg_3109_pp0_iter44_reg;
            p_read_33_reg_3109_pp0_iter46_reg <= p_read_33_reg_3109_pp0_iter45_reg;
            p_read_33_reg_3109_pp0_iter47_reg <= p_read_33_reg_3109_pp0_iter46_reg;
            p_read_33_reg_3109_pp0_iter48_reg <= p_read_33_reg_3109_pp0_iter47_reg;
            p_read_33_reg_3109_pp0_iter49_reg <= p_read_33_reg_3109_pp0_iter48_reg;
            p_read_33_reg_3109_pp0_iter4_reg <= p_read_33_reg_3109_pp0_iter3_reg;
            p_read_33_reg_3109_pp0_iter50_reg <= p_read_33_reg_3109_pp0_iter49_reg;
            p_read_33_reg_3109_pp0_iter51_reg <= p_read_33_reg_3109_pp0_iter50_reg;
            p_read_33_reg_3109_pp0_iter52_reg <= p_read_33_reg_3109_pp0_iter51_reg;
            p_read_33_reg_3109_pp0_iter53_reg <= p_read_33_reg_3109_pp0_iter52_reg;
            p_read_33_reg_3109_pp0_iter54_reg <= p_read_33_reg_3109_pp0_iter53_reg;
            p_read_33_reg_3109_pp0_iter55_reg <= p_read_33_reg_3109_pp0_iter54_reg;
            p_read_33_reg_3109_pp0_iter56_reg <= p_read_33_reg_3109_pp0_iter55_reg;
            p_read_33_reg_3109_pp0_iter57_reg <= p_read_33_reg_3109_pp0_iter56_reg;
            p_read_33_reg_3109_pp0_iter58_reg <= p_read_33_reg_3109_pp0_iter57_reg;
            p_read_33_reg_3109_pp0_iter59_reg <= p_read_33_reg_3109_pp0_iter58_reg;
            p_read_33_reg_3109_pp0_iter5_reg <= p_read_33_reg_3109_pp0_iter4_reg;
            p_read_33_reg_3109_pp0_iter60_reg <= p_read_33_reg_3109_pp0_iter59_reg;
            p_read_33_reg_3109_pp0_iter61_reg <= p_read_33_reg_3109_pp0_iter60_reg;
            p_read_33_reg_3109_pp0_iter62_reg <= p_read_33_reg_3109_pp0_iter61_reg;
            p_read_33_reg_3109_pp0_iter63_reg <= p_read_33_reg_3109_pp0_iter62_reg;
            p_read_33_reg_3109_pp0_iter64_reg <= p_read_33_reg_3109_pp0_iter63_reg;
            p_read_33_reg_3109_pp0_iter65_reg <= p_read_33_reg_3109_pp0_iter64_reg;
            p_read_33_reg_3109_pp0_iter66_reg <= p_read_33_reg_3109_pp0_iter65_reg;
            p_read_33_reg_3109_pp0_iter67_reg <= p_read_33_reg_3109_pp0_iter66_reg;
            p_read_33_reg_3109_pp0_iter68_reg <= p_read_33_reg_3109_pp0_iter67_reg;
            p_read_33_reg_3109_pp0_iter69_reg <= p_read_33_reg_3109_pp0_iter68_reg;
            p_read_33_reg_3109_pp0_iter6_reg <= p_read_33_reg_3109_pp0_iter5_reg;
            p_read_33_reg_3109_pp0_iter70_reg <= p_read_33_reg_3109_pp0_iter69_reg;
            p_read_33_reg_3109_pp0_iter71_reg <= p_read_33_reg_3109_pp0_iter70_reg;
            p_read_33_reg_3109_pp0_iter72_reg <= p_read_33_reg_3109_pp0_iter71_reg;
            p_read_33_reg_3109_pp0_iter73_reg <= p_read_33_reg_3109_pp0_iter72_reg;
            p_read_33_reg_3109_pp0_iter74_reg <= p_read_33_reg_3109_pp0_iter73_reg;
            p_read_33_reg_3109_pp0_iter75_reg <= p_read_33_reg_3109_pp0_iter74_reg;
            p_read_33_reg_3109_pp0_iter76_reg <= p_read_33_reg_3109_pp0_iter75_reg;
            p_read_33_reg_3109_pp0_iter7_reg <= p_read_33_reg_3109_pp0_iter6_reg;
            p_read_33_reg_3109_pp0_iter8_reg <= p_read_33_reg_3109_pp0_iter7_reg;
            p_read_33_reg_3109_pp0_iter9_reg <= p_read_33_reg_3109_pp0_iter8_reg;
            p_read_34_reg_3114 <= p_read30_int_reg;
            p_read_34_reg_3114_pp0_iter10_reg <= p_read_34_reg_3114_pp0_iter9_reg;
            p_read_34_reg_3114_pp0_iter11_reg <= p_read_34_reg_3114_pp0_iter10_reg;
            p_read_34_reg_3114_pp0_iter12_reg <= p_read_34_reg_3114_pp0_iter11_reg;
            p_read_34_reg_3114_pp0_iter13_reg <= p_read_34_reg_3114_pp0_iter12_reg;
            p_read_34_reg_3114_pp0_iter14_reg <= p_read_34_reg_3114_pp0_iter13_reg;
            p_read_34_reg_3114_pp0_iter15_reg <= p_read_34_reg_3114_pp0_iter14_reg;
            p_read_34_reg_3114_pp0_iter16_reg <= p_read_34_reg_3114_pp0_iter15_reg;
            p_read_34_reg_3114_pp0_iter17_reg <= p_read_34_reg_3114_pp0_iter16_reg;
            p_read_34_reg_3114_pp0_iter18_reg <= p_read_34_reg_3114_pp0_iter17_reg;
            p_read_34_reg_3114_pp0_iter19_reg <= p_read_34_reg_3114_pp0_iter18_reg;
            p_read_34_reg_3114_pp0_iter1_reg <= p_read_34_reg_3114;
            p_read_34_reg_3114_pp0_iter20_reg <= p_read_34_reg_3114_pp0_iter19_reg;
            p_read_34_reg_3114_pp0_iter21_reg <= p_read_34_reg_3114_pp0_iter20_reg;
            p_read_34_reg_3114_pp0_iter22_reg <= p_read_34_reg_3114_pp0_iter21_reg;
            p_read_34_reg_3114_pp0_iter23_reg <= p_read_34_reg_3114_pp0_iter22_reg;
            p_read_34_reg_3114_pp0_iter24_reg <= p_read_34_reg_3114_pp0_iter23_reg;
            p_read_34_reg_3114_pp0_iter25_reg <= p_read_34_reg_3114_pp0_iter24_reg;
            p_read_34_reg_3114_pp0_iter26_reg <= p_read_34_reg_3114_pp0_iter25_reg;
            p_read_34_reg_3114_pp0_iter27_reg <= p_read_34_reg_3114_pp0_iter26_reg;
            p_read_34_reg_3114_pp0_iter28_reg <= p_read_34_reg_3114_pp0_iter27_reg;
            p_read_34_reg_3114_pp0_iter29_reg <= p_read_34_reg_3114_pp0_iter28_reg;
            p_read_34_reg_3114_pp0_iter2_reg <= p_read_34_reg_3114_pp0_iter1_reg;
            p_read_34_reg_3114_pp0_iter30_reg <= p_read_34_reg_3114_pp0_iter29_reg;
            p_read_34_reg_3114_pp0_iter31_reg <= p_read_34_reg_3114_pp0_iter30_reg;
            p_read_34_reg_3114_pp0_iter32_reg <= p_read_34_reg_3114_pp0_iter31_reg;
            p_read_34_reg_3114_pp0_iter33_reg <= p_read_34_reg_3114_pp0_iter32_reg;
            p_read_34_reg_3114_pp0_iter34_reg <= p_read_34_reg_3114_pp0_iter33_reg;
            p_read_34_reg_3114_pp0_iter35_reg <= p_read_34_reg_3114_pp0_iter34_reg;
            p_read_34_reg_3114_pp0_iter36_reg <= p_read_34_reg_3114_pp0_iter35_reg;
            p_read_34_reg_3114_pp0_iter37_reg <= p_read_34_reg_3114_pp0_iter36_reg;
            p_read_34_reg_3114_pp0_iter38_reg <= p_read_34_reg_3114_pp0_iter37_reg;
            p_read_34_reg_3114_pp0_iter39_reg <= p_read_34_reg_3114_pp0_iter38_reg;
            p_read_34_reg_3114_pp0_iter3_reg <= p_read_34_reg_3114_pp0_iter2_reg;
            p_read_34_reg_3114_pp0_iter40_reg <= p_read_34_reg_3114_pp0_iter39_reg;
            p_read_34_reg_3114_pp0_iter41_reg <= p_read_34_reg_3114_pp0_iter40_reg;
            p_read_34_reg_3114_pp0_iter42_reg <= p_read_34_reg_3114_pp0_iter41_reg;
            p_read_34_reg_3114_pp0_iter43_reg <= p_read_34_reg_3114_pp0_iter42_reg;
            p_read_34_reg_3114_pp0_iter44_reg <= p_read_34_reg_3114_pp0_iter43_reg;
            p_read_34_reg_3114_pp0_iter45_reg <= p_read_34_reg_3114_pp0_iter44_reg;
            p_read_34_reg_3114_pp0_iter46_reg <= p_read_34_reg_3114_pp0_iter45_reg;
            p_read_34_reg_3114_pp0_iter47_reg <= p_read_34_reg_3114_pp0_iter46_reg;
            p_read_34_reg_3114_pp0_iter48_reg <= p_read_34_reg_3114_pp0_iter47_reg;
            p_read_34_reg_3114_pp0_iter49_reg <= p_read_34_reg_3114_pp0_iter48_reg;
            p_read_34_reg_3114_pp0_iter4_reg <= p_read_34_reg_3114_pp0_iter3_reg;
            p_read_34_reg_3114_pp0_iter50_reg <= p_read_34_reg_3114_pp0_iter49_reg;
            p_read_34_reg_3114_pp0_iter51_reg <= p_read_34_reg_3114_pp0_iter50_reg;
            p_read_34_reg_3114_pp0_iter52_reg <= p_read_34_reg_3114_pp0_iter51_reg;
            p_read_34_reg_3114_pp0_iter53_reg <= p_read_34_reg_3114_pp0_iter52_reg;
            p_read_34_reg_3114_pp0_iter54_reg <= p_read_34_reg_3114_pp0_iter53_reg;
            p_read_34_reg_3114_pp0_iter55_reg <= p_read_34_reg_3114_pp0_iter54_reg;
            p_read_34_reg_3114_pp0_iter56_reg <= p_read_34_reg_3114_pp0_iter55_reg;
            p_read_34_reg_3114_pp0_iter57_reg <= p_read_34_reg_3114_pp0_iter56_reg;
            p_read_34_reg_3114_pp0_iter58_reg <= p_read_34_reg_3114_pp0_iter57_reg;
            p_read_34_reg_3114_pp0_iter59_reg <= p_read_34_reg_3114_pp0_iter58_reg;
            p_read_34_reg_3114_pp0_iter5_reg <= p_read_34_reg_3114_pp0_iter4_reg;
            p_read_34_reg_3114_pp0_iter60_reg <= p_read_34_reg_3114_pp0_iter59_reg;
            p_read_34_reg_3114_pp0_iter61_reg <= p_read_34_reg_3114_pp0_iter60_reg;
            p_read_34_reg_3114_pp0_iter62_reg <= p_read_34_reg_3114_pp0_iter61_reg;
            p_read_34_reg_3114_pp0_iter63_reg <= p_read_34_reg_3114_pp0_iter62_reg;
            p_read_34_reg_3114_pp0_iter64_reg <= p_read_34_reg_3114_pp0_iter63_reg;
            p_read_34_reg_3114_pp0_iter65_reg <= p_read_34_reg_3114_pp0_iter64_reg;
            p_read_34_reg_3114_pp0_iter66_reg <= p_read_34_reg_3114_pp0_iter65_reg;
            p_read_34_reg_3114_pp0_iter67_reg <= p_read_34_reg_3114_pp0_iter66_reg;
            p_read_34_reg_3114_pp0_iter68_reg <= p_read_34_reg_3114_pp0_iter67_reg;
            p_read_34_reg_3114_pp0_iter69_reg <= p_read_34_reg_3114_pp0_iter68_reg;
            p_read_34_reg_3114_pp0_iter6_reg <= p_read_34_reg_3114_pp0_iter5_reg;
            p_read_34_reg_3114_pp0_iter70_reg <= p_read_34_reg_3114_pp0_iter69_reg;
            p_read_34_reg_3114_pp0_iter71_reg <= p_read_34_reg_3114_pp0_iter70_reg;
            p_read_34_reg_3114_pp0_iter72_reg <= p_read_34_reg_3114_pp0_iter71_reg;
            p_read_34_reg_3114_pp0_iter73_reg <= p_read_34_reg_3114_pp0_iter72_reg;
            p_read_34_reg_3114_pp0_iter74_reg <= p_read_34_reg_3114_pp0_iter73_reg;
            p_read_34_reg_3114_pp0_iter75_reg <= p_read_34_reg_3114_pp0_iter74_reg;
            p_read_34_reg_3114_pp0_iter76_reg <= p_read_34_reg_3114_pp0_iter75_reg;
            p_read_34_reg_3114_pp0_iter7_reg <= p_read_34_reg_3114_pp0_iter6_reg;
            p_read_34_reg_3114_pp0_iter8_reg <= p_read_34_reg_3114_pp0_iter7_reg;
            p_read_34_reg_3114_pp0_iter9_reg <= p_read_34_reg_3114_pp0_iter8_reg;
            p_read_35_reg_3119 <= p_read29_int_reg;
            p_read_35_reg_3119_pp0_iter10_reg <= p_read_35_reg_3119_pp0_iter9_reg;
            p_read_35_reg_3119_pp0_iter11_reg <= p_read_35_reg_3119_pp0_iter10_reg;
            p_read_35_reg_3119_pp0_iter12_reg <= p_read_35_reg_3119_pp0_iter11_reg;
            p_read_35_reg_3119_pp0_iter13_reg <= p_read_35_reg_3119_pp0_iter12_reg;
            p_read_35_reg_3119_pp0_iter14_reg <= p_read_35_reg_3119_pp0_iter13_reg;
            p_read_35_reg_3119_pp0_iter15_reg <= p_read_35_reg_3119_pp0_iter14_reg;
            p_read_35_reg_3119_pp0_iter16_reg <= p_read_35_reg_3119_pp0_iter15_reg;
            p_read_35_reg_3119_pp0_iter17_reg <= p_read_35_reg_3119_pp0_iter16_reg;
            p_read_35_reg_3119_pp0_iter18_reg <= p_read_35_reg_3119_pp0_iter17_reg;
            p_read_35_reg_3119_pp0_iter19_reg <= p_read_35_reg_3119_pp0_iter18_reg;
            p_read_35_reg_3119_pp0_iter1_reg <= p_read_35_reg_3119;
            p_read_35_reg_3119_pp0_iter20_reg <= p_read_35_reg_3119_pp0_iter19_reg;
            p_read_35_reg_3119_pp0_iter21_reg <= p_read_35_reg_3119_pp0_iter20_reg;
            p_read_35_reg_3119_pp0_iter22_reg <= p_read_35_reg_3119_pp0_iter21_reg;
            p_read_35_reg_3119_pp0_iter23_reg <= p_read_35_reg_3119_pp0_iter22_reg;
            p_read_35_reg_3119_pp0_iter24_reg <= p_read_35_reg_3119_pp0_iter23_reg;
            p_read_35_reg_3119_pp0_iter25_reg <= p_read_35_reg_3119_pp0_iter24_reg;
            p_read_35_reg_3119_pp0_iter26_reg <= p_read_35_reg_3119_pp0_iter25_reg;
            p_read_35_reg_3119_pp0_iter27_reg <= p_read_35_reg_3119_pp0_iter26_reg;
            p_read_35_reg_3119_pp0_iter28_reg <= p_read_35_reg_3119_pp0_iter27_reg;
            p_read_35_reg_3119_pp0_iter29_reg <= p_read_35_reg_3119_pp0_iter28_reg;
            p_read_35_reg_3119_pp0_iter2_reg <= p_read_35_reg_3119_pp0_iter1_reg;
            p_read_35_reg_3119_pp0_iter30_reg <= p_read_35_reg_3119_pp0_iter29_reg;
            p_read_35_reg_3119_pp0_iter31_reg <= p_read_35_reg_3119_pp0_iter30_reg;
            p_read_35_reg_3119_pp0_iter32_reg <= p_read_35_reg_3119_pp0_iter31_reg;
            p_read_35_reg_3119_pp0_iter33_reg <= p_read_35_reg_3119_pp0_iter32_reg;
            p_read_35_reg_3119_pp0_iter34_reg <= p_read_35_reg_3119_pp0_iter33_reg;
            p_read_35_reg_3119_pp0_iter35_reg <= p_read_35_reg_3119_pp0_iter34_reg;
            p_read_35_reg_3119_pp0_iter36_reg <= p_read_35_reg_3119_pp0_iter35_reg;
            p_read_35_reg_3119_pp0_iter37_reg <= p_read_35_reg_3119_pp0_iter36_reg;
            p_read_35_reg_3119_pp0_iter38_reg <= p_read_35_reg_3119_pp0_iter37_reg;
            p_read_35_reg_3119_pp0_iter39_reg <= p_read_35_reg_3119_pp0_iter38_reg;
            p_read_35_reg_3119_pp0_iter3_reg <= p_read_35_reg_3119_pp0_iter2_reg;
            p_read_35_reg_3119_pp0_iter40_reg <= p_read_35_reg_3119_pp0_iter39_reg;
            p_read_35_reg_3119_pp0_iter41_reg <= p_read_35_reg_3119_pp0_iter40_reg;
            p_read_35_reg_3119_pp0_iter42_reg <= p_read_35_reg_3119_pp0_iter41_reg;
            p_read_35_reg_3119_pp0_iter43_reg <= p_read_35_reg_3119_pp0_iter42_reg;
            p_read_35_reg_3119_pp0_iter44_reg <= p_read_35_reg_3119_pp0_iter43_reg;
            p_read_35_reg_3119_pp0_iter45_reg <= p_read_35_reg_3119_pp0_iter44_reg;
            p_read_35_reg_3119_pp0_iter46_reg <= p_read_35_reg_3119_pp0_iter45_reg;
            p_read_35_reg_3119_pp0_iter47_reg <= p_read_35_reg_3119_pp0_iter46_reg;
            p_read_35_reg_3119_pp0_iter48_reg <= p_read_35_reg_3119_pp0_iter47_reg;
            p_read_35_reg_3119_pp0_iter49_reg <= p_read_35_reg_3119_pp0_iter48_reg;
            p_read_35_reg_3119_pp0_iter4_reg <= p_read_35_reg_3119_pp0_iter3_reg;
            p_read_35_reg_3119_pp0_iter50_reg <= p_read_35_reg_3119_pp0_iter49_reg;
            p_read_35_reg_3119_pp0_iter51_reg <= p_read_35_reg_3119_pp0_iter50_reg;
            p_read_35_reg_3119_pp0_iter52_reg <= p_read_35_reg_3119_pp0_iter51_reg;
            p_read_35_reg_3119_pp0_iter53_reg <= p_read_35_reg_3119_pp0_iter52_reg;
            p_read_35_reg_3119_pp0_iter54_reg <= p_read_35_reg_3119_pp0_iter53_reg;
            p_read_35_reg_3119_pp0_iter55_reg <= p_read_35_reg_3119_pp0_iter54_reg;
            p_read_35_reg_3119_pp0_iter56_reg <= p_read_35_reg_3119_pp0_iter55_reg;
            p_read_35_reg_3119_pp0_iter57_reg <= p_read_35_reg_3119_pp0_iter56_reg;
            p_read_35_reg_3119_pp0_iter58_reg <= p_read_35_reg_3119_pp0_iter57_reg;
            p_read_35_reg_3119_pp0_iter59_reg <= p_read_35_reg_3119_pp0_iter58_reg;
            p_read_35_reg_3119_pp0_iter5_reg <= p_read_35_reg_3119_pp0_iter4_reg;
            p_read_35_reg_3119_pp0_iter60_reg <= p_read_35_reg_3119_pp0_iter59_reg;
            p_read_35_reg_3119_pp0_iter61_reg <= p_read_35_reg_3119_pp0_iter60_reg;
            p_read_35_reg_3119_pp0_iter62_reg <= p_read_35_reg_3119_pp0_iter61_reg;
            p_read_35_reg_3119_pp0_iter63_reg <= p_read_35_reg_3119_pp0_iter62_reg;
            p_read_35_reg_3119_pp0_iter64_reg <= p_read_35_reg_3119_pp0_iter63_reg;
            p_read_35_reg_3119_pp0_iter65_reg <= p_read_35_reg_3119_pp0_iter64_reg;
            p_read_35_reg_3119_pp0_iter66_reg <= p_read_35_reg_3119_pp0_iter65_reg;
            p_read_35_reg_3119_pp0_iter67_reg <= p_read_35_reg_3119_pp0_iter66_reg;
            p_read_35_reg_3119_pp0_iter68_reg <= p_read_35_reg_3119_pp0_iter67_reg;
            p_read_35_reg_3119_pp0_iter69_reg <= p_read_35_reg_3119_pp0_iter68_reg;
            p_read_35_reg_3119_pp0_iter6_reg <= p_read_35_reg_3119_pp0_iter5_reg;
            p_read_35_reg_3119_pp0_iter70_reg <= p_read_35_reg_3119_pp0_iter69_reg;
            p_read_35_reg_3119_pp0_iter71_reg <= p_read_35_reg_3119_pp0_iter70_reg;
            p_read_35_reg_3119_pp0_iter72_reg <= p_read_35_reg_3119_pp0_iter71_reg;
            p_read_35_reg_3119_pp0_iter73_reg <= p_read_35_reg_3119_pp0_iter72_reg;
            p_read_35_reg_3119_pp0_iter74_reg <= p_read_35_reg_3119_pp0_iter73_reg;
            p_read_35_reg_3119_pp0_iter75_reg <= p_read_35_reg_3119_pp0_iter74_reg;
            p_read_35_reg_3119_pp0_iter76_reg <= p_read_35_reg_3119_pp0_iter75_reg;
            p_read_35_reg_3119_pp0_iter7_reg <= p_read_35_reg_3119_pp0_iter6_reg;
            p_read_35_reg_3119_pp0_iter8_reg <= p_read_35_reg_3119_pp0_iter7_reg;
            p_read_35_reg_3119_pp0_iter9_reg <= p_read_35_reg_3119_pp0_iter8_reg;
            p_read_36_reg_3124 <= p_read28_int_reg;
            p_read_36_reg_3124_pp0_iter10_reg <= p_read_36_reg_3124_pp0_iter9_reg;
            p_read_36_reg_3124_pp0_iter11_reg <= p_read_36_reg_3124_pp0_iter10_reg;
            p_read_36_reg_3124_pp0_iter12_reg <= p_read_36_reg_3124_pp0_iter11_reg;
            p_read_36_reg_3124_pp0_iter13_reg <= p_read_36_reg_3124_pp0_iter12_reg;
            p_read_36_reg_3124_pp0_iter14_reg <= p_read_36_reg_3124_pp0_iter13_reg;
            p_read_36_reg_3124_pp0_iter15_reg <= p_read_36_reg_3124_pp0_iter14_reg;
            p_read_36_reg_3124_pp0_iter16_reg <= p_read_36_reg_3124_pp0_iter15_reg;
            p_read_36_reg_3124_pp0_iter17_reg <= p_read_36_reg_3124_pp0_iter16_reg;
            p_read_36_reg_3124_pp0_iter18_reg <= p_read_36_reg_3124_pp0_iter17_reg;
            p_read_36_reg_3124_pp0_iter19_reg <= p_read_36_reg_3124_pp0_iter18_reg;
            p_read_36_reg_3124_pp0_iter1_reg <= p_read_36_reg_3124;
            p_read_36_reg_3124_pp0_iter20_reg <= p_read_36_reg_3124_pp0_iter19_reg;
            p_read_36_reg_3124_pp0_iter21_reg <= p_read_36_reg_3124_pp0_iter20_reg;
            p_read_36_reg_3124_pp0_iter22_reg <= p_read_36_reg_3124_pp0_iter21_reg;
            p_read_36_reg_3124_pp0_iter23_reg <= p_read_36_reg_3124_pp0_iter22_reg;
            p_read_36_reg_3124_pp0_iter24_reg <= p_read_36_reg_3124_pp0_iter23_reg;
            p_read_36_reg_3124_pp0_iter25_reg <= p_read_36_reg_3124_pp0_iter24_reg;
            p_read_36_reg_3124_pp0_iter26_reg <= p_read_36_reg_3124_pp0_iter25_reg;
            p_read_36_reg_3124_pp0_iter27_reg <= p_read_36_reg_3124_pp0_iter26_reg;
            p_read_36_reg_3124_pp0_iter28_reg <= p_read_36_reg_3124_pp0_iter27_reg;
            p_read_36_reg_3124_pp0_iter29_reg <= p_read_36_reg_3124_pp0_iter28_reg;
            p_read_36_reg_3124_pp0_iter2_reg <= p_read_36_reg_3124_pp0_iter1_reg;
            p_read_36_reg_3124_pp0_iter30_reg <= p_read_36_reg_3124_pp0_iter29_reg;
            p_read_36_reg_3124_pp0_iter31_reg <= p_read_36_reg_3124_pp0_iter30_reg;
            p_read_36_reg_3124_pp0_iter32_reg <= p_read_36_reg_3124_pp0_iter31_reg;
            p_read_36_reg_3124_pp0_iter33_reg <= p_read_36_reg_3124_pp0_iter32_reg;
            p_read_36_reg_3124_pp0_iter34_reg <= p_read_36_reg_3124_pp0_iter33_reg;
            p_read_36_reg_3124_pp0_iter35_reg <= p_read_36_reg_3124_pp0_iter34_reg;
            p_read_36_reg_3124_pp0_iter36_reg <= p_read_36_reg_3124_pp0_iter35_reg;
            p_read_36_reg_3124_pp0_iter37_reg <= p_read_36_reg_3124_pp0_iter36_reg;
            p_read_36_reg_3124_pp0_iter38_reg <= p_read_36_reg_3124_pp0_iter37_reg;
            p_read_36_reg_3124_pp0_iter39_reg <= p_read_36_reg_3124_pp0_iter38_reg;
            p_read_36_reg_3124_pp0_iter3_reg <= p_read_36_reg_3124_pp0_iter2_reg;
            p_read_36_reg_3124_pp0_iter40_reg <= p_read_36_reg_3124_pp0_iter39_reg;
            p_read_36_reg_3124_pp0_iter41_reg <= p_read_36_reg_3124_pp0_iter40_reg;
            p_read_36_reg_3124_pp0_iter42_reg <= p_read_36_reg_3124_pp0_iter41_reg;
            p_read_36_reg_3124_pp0_iter43_reg <= p_read_36_reg_3124_pp0_iter42_reg;
            p_read_36_reg_3124_pp0_iter44_reg <= p_read_36_reg_3124_pp0_iter43_reg;
            p_read_36_reg_3124_pp0_iter45_reg <= p_read_36_reg_3124_pp0_iter44_reg;
            p_read_36_reg_3124_pp0_iter46_reg <= p_read_36_reg_3124_pp0_iter45_reg;
            p_read_36_reg_3124_pp0_iter47_reg <= p_read_36_reg_3124_pp0_iter46_reg;
            p_read_36_reg_3124_pp0_iter48_reg <= p_read_36_reg_3124_pp0_iter47_reg;
            p_read_36_reg_3124_pp0_iter49_reg <= p_read_36_reg_3124_pp0_iter48_reg;
            p_read_36_reg_3124_pp0_iter4_reg <= p_read_36_reg_3124_pp0_iter3_reg;
            p_read_36_reg_3124_pp0_iter50_reg <= p_read_36_reg_3124_pp0_iter49_reg;
            p_read_36_reg_3124_pp0_iter51_reg <= p_read_36_reg_3124_pp0_iter50_reg;
            p_read_36_reg_3124_pp0_iter52_reg <= p_read_36_reg_3124_pp0_iter51_reg;
            p_read_36_reg_3124_pp0_iter53_reg <= p_read_36_reg_3124_pp0_iter52_reg;
            p_read_36_reg_3124_pp0_iter54_reg <= p_read_36_reg_3124_pp0_iter53_reg;
            p_read_36_reg_3124_pp0_iter55_reg <= p_read_36_reg_3124_pp0_iter54_reg;
            p_read_36_reg_3124_pp0_iter56_reg <= p_read_36_reg_3124_pp0_iter55_reg;
            p_read_36_reg_3124_pp0_iter57_reg <= p_read_36_reg_3124_pp0_iter56_reg;
            p_read_36_reg_3124_pp0_iter58_reg <= p_read_36_reg_3124_pp0_iter57_reg;
            p_read_36_reg_3124_pp0_iter59_reg <= p_read_36_reg_3124_pp0_iter58_reg;
            p_read_36_reg_3124_pp0_iter5_reg <= p_read_36_reg_3124_pp0_iter4_reg;
            p_read_36_reg_3124_pp0_iter60_reg <= p_read_36_reg_3124_pp0_iter59_reg;
            p_read_36_reg_3124_pp0_iter61_reg <= p_read_36_reg_3124_pp0_iter60_reg;
            p_read_36_reg_3124_pp0_iter62_reg <= p_read_36_reg_3124_pp0_iter61_reg;
            p_read_36_reg_3124_pp0_iter63_reg <= p_read_36_reg_3124_pp0_iter62_reg;
            p_read_36_reg_3124_pp0_iter64_reg <= p_read_36_reg_3124_pp0_iter63_reg;
            p_read_36_reg_3124_pp0_iter65_reg <= p_read_36_reg_3124_pp0_iter64_reg;
            p_read_36_reg_3124_pp0_iter66_reg <= p_read_36_reg_3124_pp0_iter65_reg;
            p_read_36_reg_3124_pp0_iter67_reg <= p_read_36_reg_3124_pp0_iter66_reg;
            p_read_36_reg_3124_pp0_iter68_reg <= p_read_36_reg_3124_pp0_iter67_reg;
            p_read_36_reg_3124_pp0_iter69_reg <= p_read_36_reg_3124_pp0_iter68_reg;
            p_read_36_reg_3124_pp0_iter6_reg <= p_read_36_reg_3124_pp0_iter5_reg;
            p_read_36_reg_3124_pp0_iter70_reg <= p_read_36_reg_3124_pp0_iter69_reg;
            p_read_36_reg_3124_pp0_iter71_reg <= p_read_36_reg_3124_pp0_iter70_reg;
            p_read_36_reg_3124_pp0_iter72_reg <= p_read_36_reg_3124_pp0_iter71_reg;
            p_read_36_reg_3124_pp0_iter73_reg <= p_read_36_reg_3124_pp0_iter72_reg;
            p_read_36_reg_3124_pp0_iter74_reg <= p_read_36_reg_3124_pp0_iter73_reg;
            p_read_36_reg_3124_pp0_iter75_reg <= p_read_36_reg_3124_pp0_iter74_reg;
            p_read_36_reg_3124_pp0_iter76_reg <= p_read_36_reg_3124_pp0_iter75_reg;
            p_read_36_reg_3124_pp0_iter7_reg <= p_read_36_reg_3124_pp0_iter6_reg;
            p_read_36_reg_3124_pp0_iter8_reg <= p_read_36_reg_3124_pp0_iter7_reg;
            p_read_36_reg_3124_pp0_iter9_reg <= p_read_36_reg_3124_pp0_iter8_reg;
            p_read_37_reg_3129 <= p_read27_int_reg;
            p_read_37_reg_3129_pp0_iter10_reg <= p_read_37_reg_3129_pp0_iter9_reg;
            p_read_37_reg_3129_pp0_iter11_reg <= p_read_37_reg_3129_pp0_iter10_reg;
            p_read_37_reg_3129_pp0_iter12_reg <= p_read_37_reg_3129_pp0_iter11_reg;
            p_read_37_reg_3129_pp0_iter13_reg <= p_read_37_reg_3129_pp0_iter12_reg;
            p_read_37_reg_3129_pp0_iter14_reg <= p_read_37_reg_3129_pp0_iter13_reg;
            p_read_37_reg_3129_pp0_iter15_reg <= p_read_37_reg_3129_pp0_iter14_reg;
            p_read_37_reg_3129_pp0_iter16_reg <= p_read_37_reg_3129_pp0_iter15_reg;
            p_read_37_reg_3129_pp0_iter17_reg <= p_read_37_reg_3129_pp0_iter16_reg;
            p_read_37_reg_3129_pp0_iter18_reg <= p_read_37_reg_3129_pp0_iter17_reg;
            p_read_37_reg_3129_pp0_iter19_reg <= p_read_37_reg_3129_pp0_iter18_reg;
            p_read_37_reg_3129_pp0_iter1_reg <= p_read_37_reg_3129;
            p_read_37_reg_3129_pp0_iter20_reg <= p_read_37_reg_3129_pp0_iter19_reg;
            p_read_37_reg_3129_pp0_iter21_reg <= p_read_37_reg_3129_pp0_iter20_reg;
            p_read_37_reg_3129_pp0_iter22_reg <= p_read_37_reg_3129_pp0_iter21_reg;
            p_read_37_reg_3129_pp0_iter23_reg <= p_read_37_reg_3129_pp0_iter22_reg;
            p_read_37_reg_3129_pp0_iter24_reg <= p_read_37_reg_3129_pp0_iter23_reg;
            p_read_37_reg_3129_pp0_iter25_reg <= p_read_37_reg_3129_pp0_iter24_reg;
            p_read_37_reg_3129_pp0_iter26_reg <= p_read_37_reg_3129_pp0_iter25_reg;
            p_read_37_reg_3129_pp0_iter27_reg <= p_read_37_reg_3129_pp0_iter26_reg;
            p_read_37_reg_3129_pp0_iter28_reg <= p_read_37_reg_3129_pp0_iter27_reg;
            p_read_37_reg_3129_pp0_iter29_reg <= p_read_37_reg_3129_pp0_iter28_reg;
            p_read_37_reg_3129_pp0_iter2_reg <= p_read_37_reg_3129_pp0_iter1_reg;
            p_read_37_reg_3129_pp0_iter30_reg <= p_read_37_reg_3129_pp0_iter29_reg;
            p_read_37_reg_3129_pp0_iter31_reg <= p_read_37_reg_3129_pp0_iter30_reg;
            p_read_37_reg_3129_pp0_iter32_reg <= p_read_37_reg_3129_pp0_iter31_reg;
            p_read_37_reg_3129_pp0_iter33_reg <= p_read_37_reg_3129_pp0_iter32_reg;
            p_read_37_reg_3129_pp0_iter34_reg <= p_read_37_reg_3129_pp0_iter33_reg;
            p_read_37_reg_3129_pp0_iter35_reg <= p_read_37_reg_3129_pp0_iter34_reg;
            p_read_37_reg_3129_pp0_iter36_reg <= p_read_37_reg_3129_pp0_iter35_reg;
            p_read_37_reg_3129_pp0_iter37_reg <= p_read_37_reg_3129_pp0_iter36_reg;
            p_read_37_reg_3129_pp0_iter38_reg <= p_read_37_reg_3129_pp0_iter37_reg;
            p_read_37_reg_3129_pp0_iter39_reg <= p_read_37_reg_3129_pp0_iter38_reg;
            p_read_37_reg_3129_pp0_iter3_reg <= p_read_37_reg_3129_pp0_iter2_reg;
            p_read_37_reg_3129_pp0_iter40_reg <= p_read_37_reg_3129_pp0_iter39_reg;
            p_read_37_reg_3129_pp0_iter41_reg <= p_read_37_reg_3129_pp0_iter40_reg;
            p_read_37_reg_3129_pp0_iter42_reg <= p_read_37_reg_3129_pp0_iter41_reg;
            p_read_37_reg_3129_pp0_iter43_reg <= p_read_37_reg_3129_pp0_iter42_reg;
            p_read_37_reg_3129_pp0_iter44_reg <= p_read_37_reg_3129_pp0_iter43_reg;
            p_read_37_reg_3129_pp0_iter45_reg <= p_read_37_reg_3129_pp0_iter44_reg;
            p_read_37_reg_3129_pp0_iter46_reg <= p_read_37_reg_3129_pp0_iter45_reg;
            p_read_37_reg_3129_pp0_iter47_reg <= p_read_37_reg_3129_pp0_iter46_reg;
            p_read_37_reg_3129_pp0_iter48_reg <= p_read_37_reg_3129_pp0_iter47_reg;
            p_read_37_reg_3129_pp0_iter49_reg <= p_read_37_reg_3129_pp0_iter48_reg;
            p_read_37_reg_3129_pp0_iter4_reg <= p_read_37_reg_3129_pp0_iter3_reg;
            p_read_37_reg_3129_pp0_iter50_reg <= p_read_37_reg_3129_pp0_iter49_reg;
            p_read_37_reg_3129_pp0_iter51_reg <= p_read_37_reg_3129_pp0_iter50_reg;
            p_read_37_reg_3129_pp0_iter52_reg <= p_read_37_reg_3129_pp0_iter51_reg;
            p_read_37_reg_3129_pp0_iter53_reg <= p_read_37_reg_3129_pp0_iter52_reg;
            p_read_37_reg_3129_pp0_iter54_reg <= p_read_37_reg_3129_pp0_iter53_reg;
            p_read_37_reg_3129_pp0_iter55_reg <= p_read_37_reg_3129_pp0_iter54_reg;
            p_read_37_reg_3129_pp0_iter56_reg <= p_read_37_reg_3129_pp0_iter55_reg;
            p_read_37_reg_3129_pp0_iter57_reg <= p_read_37_reg_3129_pp0_iter56_reg;
            p_read_37_reg_3129_pp0_iter58_reg <= p_read_37_reg_3129_pp0_iter57_reg;
            p_read_37_reg_3129_pp0_iter59_reg <= p_read_37_reg_3129_pp0_iter58_reg;
            p_read_37_reg_3129_pp0_iter5_reg <= p_read_37_reg_3129_pp0_iter4_reg;
            p_read_37_reg_3129_pp0_iter60_reg <= p_read_37_reg_3129_pp0_iter59_reg;
            p_read_37_reg_3129_pp0_iter61_reg <= p_read_37_reg_3129_pp0_iter60_reg;
            p_read_37_reg_3129_pp0_iter62_reg <= p_read_37_reg_3129_pp0_iter61_reg;
            p_read_37_reg_3129_pp0_iter63_reg <= p_read_37_reg_3129_pp0_iter62_reg;
            p_read_37_reg_3129_pp0_iter64_reg <= p_read_37_reg_3129_pp0_iter63_reg;
            p_read_37_reg_3129_pp0_iter65_reg <= p_read_37_reg_3129_pp0_iter64_reg;
            p_read_37_reg_3129_pp0_iter66_reg <= p_read_37_reg_3129_pp0_iter65_reg;
            p_read_37_reg_3129_pp0_iter67_reg <= p_read_37_reg_3129_pp0_iter66_reg;
            p_read_37_reg_3129_pp0_iter68_reg <= p_read_37_reg_3129_pp0_iter67_reg;
            p_read_37_reg_3129_pp0_iter69_reg <= p_read_37_reg_3129_pp0_iter68_reg;
            p_read_37_reg_3129_pp0_iter6_reg <= p_read_37_reg_3129_pp0_iter5_reg;
            p_read_37_reg_3129_pp0_iter70_reg <= p_read_37_reg_3129_pp0_iter69_reg;
            p_read_37_reg_3129_pp0_iter71_reg <= p_read_37_reg_3129_pp0_iter70_reg;
            p_read_37_reg_3129_pp0_iter72_reg <= p_read_37_reg_3129_pp0_iter71_reg;
            p_read_37_reg_3129_pp0_iter73_reg <= p_read_37_reg_3129_pp0_iter72_reg;
            p_read_37_reg_3129_pp0_iter74_reg <= p_read_37_reg_3129_pp0_iter73_reg;
            p_read_37_reg_3129_pp0_iter75_reg <= p_read_37_reg_3129_pp0_iter74_reg;
            p_read_37_reg_3129_pp0_iter76_reg <= p_read_37_reg_3129_pp0_iter75_reg;
            p_read_37_reg_3129_pp0_iter7_reg <= p_read_37_reg_3129_pp0_iter6_reg;
            p_read_37_reg_3129_pp0_iter8_reg <= p_read_37_reg_3129_pp0_iter7_reg;
            p_read_37_reg_3129_pp0_iter9_reg <= p_read_37_reg_3129_pp0_iter8_reg;
            p_read_38_reg_3134 <= p_read26_int_reg;
            p_read_38_reg_3134_pp0_iter10_reg <= p_read_38_reg_3134_pp0_iter9_reg;
            p_read_38_reg_3134_pp0_iter11_reg <= p_read_38_reg_3134_pp0_iter10_reg;
            p_read_38_reg_3134_pp0_iter12_reg <= p_read_38_reg_3134_pp0_iter11_reg;
            p_read_38_reg_3134_pp0_iter13_reg <= p_read_38_reg_3134_pp0_iter12_reg;
            p_read_38_reg_3134_pp0_iter14_reg <= p_read_38_reg_3134_pp0_iter13_reg;
            p_read_38_reg_3134_pp0_iter15_reg <= p_read_38_reg_3134_pp0_iter14_reg;
            p_read_38_reg_3134_pp0_iter16_reg <= p_read_38_reg_3134_pp0_iter15_reg;
            p_read_38_reg_3134_pp0_iter17_reg <= p_read_38_reg_3134_pp0_iter16_reg;
            p_read_38_reg_3134_pp0_iter18_reg <= p_read_38_reg_3134_pp0_iter17_reg;
            p_read_38_reg_3134_pp0_iter19_reg <= p_read_38_reg_3134_pp0_iter18_reg;
            p_read_38_reg_3134_pp0_iter1_reg <= p_read_38_reg_3134;
            p_read_38_reg_3134_pp0_iter20_reg <= p_read_38_reg_3134_pp0_iter19_reg;
            p_read_38_reg_3134_pp0_iter21_reg <= p_read_38_reg_3134_pp0_iter20_reg;
            p_read_38_reg_3134_pp0_iter22_reg <= p_read_38_reg_3134_pp0_iter21_reg;
            p_read_38_reg_3134_pp0_iter23_reg <= p_read_38_reg_3134_pp0_iter22_reg;
            p_read_38_reg_3134_pp0_iter24_reg <= p_read_38_reg_3134_pp0_iter23_reg;
            p_read_38_reg_3134_pp0_iter25_reg <= p_read_38_reg_3134_pp0_iter24_reg;
            p_read_38_reg_3134_pp0_iter26_reg <= p_read_38_reg_3134_pp0_iter25_reg;
            p_read_38_reg_3134_pp0_iter27_reg <= p_read_38_reg_3134_pp0_iter26_reg;
            p_read_38_reg_3134_pp0_iter28_reg <= p_read_38_reg_3134_pp0_iter27_reg;
            p_read_38_reg_3134_pp0_iter29_reg <= p_read_38_reg_3134_pp0_iter28_reg;
            p_read_38_reg_3134_pp0_iter2_reg <= p_read_38_reg_3134_pp0_iter1_reg;
            p_read_38_reg_3134_pp0_iter30_reg <= p_read_38_reg_3134_pp0_iter29_reg;
            p_read_38_reg_3134_pp0_iter31_reg <= p_read_38_reg_3134_pp0_iter30_reg;
            p_read_38_reg_3134_pp0_iter32_reg <= p_read_38_reg_3134_pp0_iter31_reg;
            p_read_38_reg_3134_pp0_iter33_reg <= p_read_38_reg_3134_pp0_iter32_reg;
            p_read_38_reg_3134_pp0_iter34_reg <= p_read_38_reg_3134_pp0_iter33_reg;
            p_read_38_reg_3134_pp0_iter35_reg <= p_read_38_reg_3134_pp0_iter34_reg;
            p_read_38_reg_3134_pp0_iter36_reg <= p_read_38_reg_3134_pp0_iter35_reg;
            p_read_38_reg_3134_pp0_iter37_reg <= p_read_38_reg_3134_pp0_iter36_reg;
            p_read_38_reg_3134_pp0_iter38_reg <= p_read_38_reg_3134_pp0_iter37_reg;
            p_read_38_reg_3134_pp0_iter39_reg <= p_read_38_reg_3134_pp0_iter38_reg;
            p_read_38_reg_3134_pp0_iter3_reg <= p_read_38_reg_3134_pp0_iter2_reg;
            p_read_38_reg_3134_pp0_iter40_reg <= p_read_38_reg_3134_pp0_iter39_reg;
            p_read_38_reg_3134_pp0_iter41_reg <= p_read_38_reg_3134_pp0_iter40_reg;
            p_read_38_reg_3134_pp0_iter42_reg <= p_read_38_reg_3134_pp0_iter41_reg;
            p_read_38_reg_3134_pp0_iter43_reg <= p_read_38_reg_3134_pp0_iter42_reg;
            p_read_38_reg_3134_pp0_iter44_reg <= p_read_38_reg_3134_pp0_iter43_reg;
            p_read_38_reg_3134_pp0_iter45_reg <= p_read_38_reg_3134_pp0_iter44_reg;
            p_read_38_reg_3134_pp0_iter46_reg <= p_read_38_reg_3134_pp0_iter45_reg;
            p_read_38_reg_3134_pp0_iter47_reg <= p_read_38_reg_3134_pp0_iter46_reg;
            p_read_38_reg_3134_pp0_iter48_reg <= p_read_38_reg_3134_pp0_iter47_reg;
            p_read_38_reg_3134_pp0_iter49_reg <= p_read_38_reg_3134_pp0_iter48_reg;
            p_read_38_reg_3134_pp0_iter4_reg <= p_read_38_reg_3134_pp0_iter3_reg;
            p_read_38_reg_3134_pp0_iter50_reg <= p_read_38_reg_3134_pp0_iter49_reg;
            p_read_38_reg_3134_pp0_iter51_reg <= p_read_38_reg_3134_pp0_iter50_reg;
            p_read_38_reg_3134_pp0_iter52_reg <= p_read_38_reg_3134_pp0_iter51_reg;
            p_read_38_reg_3134_pp0_iter53_reg <= p_read_38_reg_3134_pp0_iter52_reg;
            p_read_38_reg_3134_pp0_iter54_reg <= p_read_38_reg_3134_pp0_iter53_reg;
            p_read_38_reg_3134_pp0_iter55_reg <= p_read_38_reg_3134_pp0_iter54_reg;
            p_read_38_reg_3134_pp0_iter56_reg <= p_read_38_reg_3134_pp0_iter55_reg;
            p_read_38_reg_3134_pp0_iter57_reg <= p_read_38_reg_3134_pp0_iter56_reg;
            p_read_38_reg_3134_pp0_iter58_reg <= p_read_38_reg_3134_pp0_iter57_reg;
            p_read_38_reg_3134_pp0_iter59_reg <= p_read_38_reg_3134_pp0_iter58_reg;
            p_read_38_reg_3134_pp0_iter5_reg <= p_read_38_reg_3134_pp0_iter4_reg;
            p_read_38_reg_3134_pp0_iter60_reg <= p_read_38_reg_3134_pp0_iter59_reg;
            p_read_38_reg_3134_pp0_iter61_reg <= p_read_38_reg_3134_pp0_iter60_reg;
            p_read_38_reg_3134_pp0_iter62_reg <= p_read_38_reg_3134_pp0_iter61_reg;
            p_read_38_reg_3134_pp0_iter63_reg <= p_read_38_reg_3134_pp0_iter62_reg;
            p_read_38_reg_3134_pp0_iter64_reg <= p_read_38_reg_3134_pp0_iter63_reg;
            p_read_38_reg_3134_pp0_iter65_reg <= p_read_38_reg_3134_pp0_iter64_reg;
            p_read_38_reg_3134_pp0_iter66_reg <= p_read_38_reg_3134_pp0_iter65_reg;
            p_read_38_reg_3134_pp0_iter67_reg <= p_read_38_reg_3134_pp0_iter66_reg;
            p_read_38_reg_3134_pp0_iter68_reg <= p_read_38_reg_3134_pp0_iter67_reg;
            p_read_38_reg_3134_pp0_iter69_reg <= p_read_38_reg_3134_pp0_iter68_reg;
            p_read_38_reg_3134_pp0_iter6_reg <= p_read_38_reg_3134_pp0_iter5_reg;
            p_read_38_reg_3134_pp0_iter70_reg <= p_read_38_reg_3134_pp0_iter69_reg;
            p_read_38_reg_3134_pp0_iter71_reg <= p_read_38_reg_3134_pp0_iter70_reg;
            p_read_38_reg_3134_pp0_iter72_reg <= p_read_38_reg_3134_pp0_iter71_reg;
            p_read_38_reg_3134_pp0_iter73_reg <= p_read_38_reg_3134_pp0_iter72_reg;
            p_read_38_reg_3134_pp0_iter74_reg <= p_read_38_reg_3134_pp0_iter73_reg;
            p_read_38_reg_3134_pp0_iter75_reg <= p_read_38_reg_3134_pp0_iter74_reg;
            p_read_38_reg_3134_pp0_iter76_reg <= p_read_38_reg_3134_pp0_iter75_reg;
            p_read_38_reg_3134_pp0_iter7_reg <= p_read_38_reg_3134_pp0_iter6_reg;
            p_read_38_reg_3134_pp0_iter8_reg <= p_read_38_reg_3134_pp0_iter7_reg;
            p_read_38_reg_3134_pp0_iter9_reg <= p_read_38_reg_3134_pp0_iter8_reg;
            p_read_39_reg_3139 <= p_read25_int_reg;
            p_read_39_reg_3139_pp0_iter10_reg <= p_read_39_reg_3139_pp0_iter9_reg;
            p_read_39_reg_3139_pp0_iter11_reg <= p_read_39_reg_3139_pp0_iter10_reg;
            p_read_39_reg_3139_pp0_iter12_reg <= p_read_39_reg_3139_pp0_iter11_reg;
            p_read_39_reg_3139_pp0_iter13_reg <= p_read_39_reg_3139_pp0_iter12_reg;
            p_read_39_reg_3139_pp0_iter14_reg <= p_read_39_reg_3139_pp0_iter13_reg;
            p_read_39_reg_3139_pp0_iter15_reg <= p_read_39_reg_3139_pp0_iter14_reg;
            p_read_39_reg_3139_pp0_iter16_reg <= p_read_39_reg_3139_pp0_iter15_reg;
            p_read_39_reg_3139_pp0_iter17_reg <= p_read_39_reg_3139_pp0_iter16_reg;
            p_read_39_reg_3139_pp0_iter18_reg <= p_read_39_reg_3139_pp0_iter17_reg;
            p_read_39_reg_3139_pp0_iter19_reg <= p_read_39_reg_3139_pp0_iter18_reg;
            p_read_39_reg_3139_pp0_iter1_reg <= p_read_39_reg_3139;
            p_read_39_reg_3139_pp0_iter20_reg <= p_read_39_reg_3139_pp0_iter19_reg;
            p_read_39_reg_3139_pp0_iter21_reg <= p_read_39_reg_3139_pp0_iter20_reg;
            p_read_39_reg_3139_pp0_iter22_reg <= p_read_39_reg_3139_pp0_iter21_reg;
            p_read_39_reg_3139_pp0_iter23_reg <= p_read_39_reg_3139_pp0_iter22_reg;
            p_read_39_reg_3139_pp0_iter24_reg <= p_read_39_reg_3139_pp0_iter23_reg;
            p_read_39_reg_3139_pp0_iter25_reg <= p_read_39_reg_3139_pp0_iter24_reg;
            p_read_39_reg_3139_pp0_iter26_reg <= p_read_39_reg_3139_pp0_iter25_reg;
            p_read_39_reg_3139_pp0_iter27_reg <= p_read_39_reg_3139_pp0_iter26_reg;
            p_read_39_reg_3139_pp0_iter28_reg <= p_read_39_reg_3139_pp0_iter27_reg;
            p_read_39_reg_3139_pp0_iter29_reg <= p_read_39_reg_3139_pp0_iter28_reg;
            p_read_39_reg_3139_pp0_iter2_reg <= p_read_39_reg_3139_pp0_iter1_reg;
            p_read_39_reg_3139_pp0_iter30_reg <= p_read_39_reg_3139_pp0_iter29_reg;
            p_read_39_reg_3139_pp0_iter31_reg <= p_read_39_reg_3139_pp0_iter30_reg;
            p_read_39_reg_3139_pp0_iter32_reg <= p_read_39_reg_3139_pp0_iter31_reg;
            p_read_39_reg_3139_pp0_iter33_reg <= p_read_39_reg_3139_pp0_iter32_reg;
            p_read_39_reg_3139_pp0_iter34_reg <= p_read_39_reg_3139_pp0_iter33_reg;
            p_read_39_reg_3139_pp0_iter35_reg <= p_read_39_reg_3139_pp0_iter34_reg;
            p_read_39_reg_3139_pp0_iter36_reg <= p_read_39_reg_3139_pp0_iter35_reg;
            p_read_39_reg_3139_pp0_iter37_reg <= p_read_39_reg_3139_pp0_iter36_reg;
            p_read_39_reg_3139_pp0_iter38_reg <= p_read_39_reg_3139_pp0_iter37_reg;
            p_read_39_reg_3139_pp0_iter39_reg <= p_read_39_reg_3139_pp0_iter38_reg;
            p_read_39_reg_3139_pp0_iter3_reg <= p_read_39_reg_3139_pp0_iter2_reg;
            p_read_39_reg_3139_pp0_iter40_reg <= p_read_39_reg_3139_pp0_iter39_reg;
            p_read_39_reg_3139_pp0_iter41_reg <= p_read_39_reg_3139_pp0_iter40_reg;
            p_read_39_reg_3139_pp0_iter42_reg <= p_read_39_reg_3139_pp0_iter41_reg;
            p_read_39_reg_3139_pp0_iter43_reg <= p_read_39_reg_3139_pp0_iter42_reg;
            p_read_39_reg_3139_pp0_iter44_reg <= p_read_39_reg_3139_pp0_iter43_reg;
            p_read_39_reg_3139_pp0_iter45_reg <= p_read_39_reg_3139_pp0_iter44_reg;
            p_read_39_reg_3139_pp0_iter46_reg <= p_read_39_reg_3139_pp0_iter45_reg;
            p_read_39_reg_3139_pp0_iter47_reg <= p_read_39_reg_3139_pp0_iter46_reg;
            p_read_39_reg_3139_pp0_iter48_reg <= p_read_39_reg_3139_pp0_iter47_reg;
            p_read_39_reg_3139_pp0_iter49_reg <= p_read_39_reg_3139_pp0_iter48_reg;
            p_read_39_reg_3139_pp0_iter4_reg <= p_read_39_reg_3139_pp0_iter3_reg;
            p_read_39_reg_3139_pp0_iter50_reg <= p_read_39_reg_3139_pp0_iter49_reg;
            p_read_39_reg_3139_pp0_iter51_reg <= p_read_39_reg_3139_pp0_iter50_reg;
            p_read_39_reg_3139_pp0_iter52_reg <= p_read_39_reg_3139_pp0_iter51_reg;
            p_read_39_reg_3139_pp0_iter53_reg <= p_read_39_reg_3139_pp0_iter52_reg;
            p_read_39_reg_3139_pp0_iter54_reg <= p_read_39_reg_3139_pp0_iter53_reg;
            p_read_39_reg_3139_pp0_iter55_reg <= p_read_39_reg_3139_pp0_iter54_reg;
            p_read_39_reg_3139_pp0_iter56_reg <= p_read_39_reg_3139_pp0_iter55_reg;
            p_read_39_reg_3139_pp0_iter57_reg <= p_read_39_reg_3139_pp0_iter56_reg;
            p_read_39_reg_3139_pp0_iter58_reg <= p_read_39_reg_3139_pp0_iter57_reg;
            p_read_39_reg_3139_pp0_iter59_reg <= p_read_39_reg_3139_pp0_iter58_reg;
            p_read_39_reg_3139_pp0_iter5_reg <= p_read_39_reg_3139_pp0_iter4_reg;
            p_read_39_reg_3139_pp0_iter60_reg <= p_read_39_reg_3139_pp0_iter59_reg;
            p_read_39_reg_3139_pp0_iter61_reg <= p_read_39_reg_3139_pp0_iter60_reg;
            p_read_39_reg_3139_pp0_iter62_reg <= p_read_39_reg_3139_pp0_iter61_reg;
            p_read_39_reg_3139_pp0_iter63_reg <= p_read_39_reg_3139_pp0_iter62_reg;
            p_read_39_reg_3139_pp0_iter64_reg <= p_read_39_reg_3139_pp0_iter63_reg;
            p_read_39_reg_3139_pp0_iter65_reg <= p_read_39_reg_3139_pp0_iter64_reg;
            p_read_39_reg_3139_pp0_iter66_reg <= p_read_39_reg_3139_pp0_iter65_reg;
            p_read_39_reg_3139_pp0_iter67_reg <= p_read_39_reg_3139_pp0_iter66_reg;
            p_read_39_reg_3139_pp0_iter68_reg <= p_read_39_reg_3139_pp0_iter67_reg;
            p_read_39_reg_3139_pp0_iter69_reg <= p_read_39_reg_3139_pp0_iter68_reg;
            p_read_39_reg_3139_pp0_iter6_reg <= p_read_39_reg_3139_pp0_iter5_reg;
            p_read_39_reg_3139_pp0_iter70_reg <= p_read_39_reg_3139_pp0_iter69_reg;
            p_read_39_reg_3139_pp0_iter71_reg <= p_read_39_reg_3139_pp0_iter70_reg;
            p_read_39_reg_3139_pp0_iter72_reg <= p_read_39_reg_3139_pp0_iter71_reg;
            p_read_39_reg_3139_pp0_iter73_reg <= p_read_39_reg_3139_pp0_iter72_reg;
            p_read_39_reg_3139_pp0_iter74_reg <= p_read_39_reg_3139_pp0_iter73_reg;
            p_read_39_reg_3139_pp0_iter75_reg <= p_read_39_reg_3139_pp0_iter74_reg;
            p_read_39_reg_3139_pp0_iter76_reg <= p_read_39_reg_3139_pp0_iter75_reg;
            p_read_39_reg_3139_pp0_iter7_reg <= p_read_39_reg_3139_pp0_iter6_reg;
            p_read_39_reg_3139_pp0_iter8_reg <= p_read_39_reg_3139_pp0_iter7_reg;
            p_read_39_reg_3139_pp0_iter9_reg <= p_read_39_reg_3139_pp0_iter8_reg;
            p_read_40_reg_3144 <= p_read24_int_reg;
            p_read_40_reg_3144_pp0_iter10_reg <= p_read_40_reg_3144_pp0_iter9_reg;
            p_read_40_reg_3144_pp0_iter11_reg <= p_read_40_reg_3144_pp0_iter10_reg;
            p_read_40_reg_3144_pp0_iter12_reg <= p_read_40_reg_3144_pp0_iter11_reg;
            p_read_40_reg_3144_pp0_iter13_reg <= p_read_40_reg_3144_pp0_iter12_reg;
            p_read_40_reg_3144_pp0_iter14_reg <= p_read_40_reg_3144_pp0_iter13_reg;
            p_read_40_reg_3144_pp0_iter15_reg <= p_read_40_reg_3144_pp0_iter14_reg;
            p_read_40_reg_3144_pp0_iter16_reg <= p_read_40_reg_3144_pp0_iter15_reg;
            p_read_40_reg_3144_pp0_iter17_reg <= p_read_40_reg_3144_pp0_iter16_reg;
            p_read_40_reg_3144_pp0_iter18_reg <= p_read_40_reg_3144_pp0_iter17_reg;
            p_read_40_reg_3144_pp0_iter19_reg <= p_read_40_reg_3144_pp0_iter18_reg;
            p_read_40_reg_3144_pp0_iter1_reg <= p_read_40_reg_3144;
            p_read_40_reg_3144_pp0_iter20_reg <= p_read_40_reg_3144_pp0_iter19_reg;
            p_read_40_reg_3144_pp0_iter21_reg <= p_read_40_reg_3144_pp0_iter20_reg;
            p_read_40_reg_3144_pp0_iter22_reg <= p_read_40_reg_3144_pp0_iter21_reg;
            p_read_40_reg_3144_pp0_iter23_reg <= p_read_40_reg_3144_pp0_iter22_reg;
            p_read_40_reg_3144_pp0_iter24_reg <= p_read_40_reg_3144_pp0_iter23_reg;
            p_read_40_reg_3144_pp0_iter25_reg <= p_read_40_reg_3144_pp0_iter24_reg;
            p_read_40_reg_3144_pp0_iter26_reg <= p_read_40_reg_3144_pp0_iter25_reg;
            p_read_40_reg_3144_pp0_iter27_reg <= p_read_40_reg_3144_pp0_iter26_reg;
            p_read_40_reg_3144_pp0_iter28_reg <= p_read_40_reg_3144_pp0_iter27_reg;
            p_read_40_reg_3144_pp0_iter29_reg <= p_read_40_reg_3144_pp0_iter28_reg;
            p_read_40_reg_3144_pp0_iter2_reg <= p_read_40_reg_3144_pp0_iter1_reg;
            p_read_40_reg_3144_pp0_iter30_reg <= p_read_40_reg_3144_pp0_iter29_reg;
            p_read_40_reg_3144_pp0_iter31_reg <= p_read_40_reg_3144_pp0_iter30_reg;
            p_read_40_reg_3144_pp0_iter32_reg <= p_read_40_reg_3144_pp0_iter31_reg;
            p_read_40_reg_3144_pp0_iter33_reg <= p_read_40_reg_3144_pp0_iter32_reg;
            p_read_40_reg_3144_pp0_iter34_reg <= p_read_40_reg_3144_pp0_iter33_reg;
            p_read_40_reg_3144_pp0_iter35_reg <= p_read_40_reg_3144_pp0_iter34_reg;
            p_read_40_reg_3144_pp0_iter36_reg <= p_read_40_reg_3144_pp0_iter35_reg;
            p_read_40_reg_3144_pp0_iter37_reg <= p_read_40_reg_3144_pp0_iter36_reg;
            p_read_40_reg_3144_pp0_iter38_reg <= p_read_40_reg_3144_pp0_iter37_reg;
            p_read_40_reg_3144_pp0_iter39_reg <= p_read_40_reg_3144_pp0_iter38_reg;
            p_read_40_reg_3144_pp0_iter3_reg <= p_read_40_reg_3144_pp0_iter2_reg;
            p_read_40_reg_3144_pp0_iter40_reg <= p_read_40_reg_3144_pp0_iter39_reg;
            p_read_40_reg_3144_pp0_iter41_reg <= p_read_40_reg_3144_pp0_iter40_reg;
            p_read_40_reg_3144_pp0_iter42_reg <= p_read_40_reg_3144_pp0_iter41_reg;
            p_read_40_reg_3144_pp0_iter43_reg <= p_read_40_reg_3144_pp0_iter42_reg;
            p_read_40_reg_3144_pp0_iter44_reg <= p_read_40_reg_3144_pp0_iter43_reg;
            p_read_40_reg_3144_pp0_iter45_reg <= p_read_40_reg_3144_pp0_iter44_reg;
            p_read_40_reg_3144_pp0_iter46_reg <= p_read_40_reg_3144_pp0_iter45_reg;
            p_read_40_reg_3144_pp0_iter47_reg <= p_read_40_reg_3144_pp0_iter46_reg;
            p_read_40_reg_3144_pp0_iter48_reg <= p_read_40_reg_3144_pp0_iter47_reg;
            p_read_40_reg_3144_pp0_iter49_reg <= p_read_40_reg_3144_pp0_iter48_reg;
            p_read_40_reg_3144_pp0_iter4_reg <= p_read_40_reg_3144_pp0_iter3_reg;
            p_read_40_reg_3144_pp0_iter50_reg <= p_read_40_reg_3144_pp0_iter49_reg;
            p_read_40_reg_3144_pp0_iter51_reg <= p_read_40_reg_3144_pp0_iter50_reg;
            p_read_40_reg_3144_pp0_iter52_reg <= p_read_40_reg_3144_pp0_iter51_reg;
            p_read_40_reg_3144_pp0_iter53_reg <= p_read_40_reg_3144_pp0_iter52_reg;
            p_read_40_reg_3144_pp0_iter54_reg <= p_read_40_reg_3144_pp0_iter53_reg;
            p_read_40_reg_3144_pp0_iter55_reg <= p_read_40_reg_3144_pp0_iter54_reg;
            p_read_40_reg_3144_pp0_iter56_reg <= p_read_40_reg_3144_pp0_iter55_reg;
            p_read_40_reg_3144_pp0_iter57_reg <= p_read_40_reg_3144_pp0_iter56_reg;
            p_read_40_reg_3144_pp0_iter58_reg <= p_read_40_reg_3144_pp0_iter57_reg;
            p_read_40_reg_3144_pp0_iter59_reg <= p_read_40_reg_3144_pp0_iter58_reg;
            p_read_40_reg_3144_pp0_iter5_reg <= p_read_40_reg_3144_pp0_iter4_reg;
            p_read_40_reg_3144_pp0_iter60_reg <= p_read_40_reg_3144_pp0_iter59_reg;
            p_read_40_reg_3144_pp0_iter61_reg <= p_read_40_reg_3144_pp0_iter60_reg;
            p_read_40_reg_3144_pp0_iter62_reg <= p_read_40_reg_3144_pp0_iter61_reg;
            p_read_40_reg_3144_pp0_iter63_reg <= p_read_40_reg_3144_pp0_iter62_reg;
            p_read_40_reg_3144_pp0_iter64_reg <= p_read_40_reg_3144_pp0_iter63_reg;
            p_read_40_reg_3144_pp0_iter65_reg <= p_read_40_reg_3144_pp0_iter64_reg;
            p_read_40_reg_3144_pp0_iter66_reg <= p_read_40_reg_3144_pp0_iter65_reg;
            p_read_40_reg_3144_pp0_iter67_reg <= p_read_40_reg_3144_pp0_iter66_reg;
            p_read_40_reg_3144_pp0_iter68_reg <= p_read_40_reg_3144_pp0_iter67_reg;
            p_read_40_reg_3144_pp0_iter69_reg <= p_read_40_reg_3144_pp0_iter68_reg;
            p_read_40_reg_3144_pp0_iter6_reg <= p_read_40_reg_3144_pp0_iter5_reg;
            p_read_40_reg_3144_pp0_iter70_reg <= p_read_40_reg_3144_pp0_iter69_reg;
            p_read_40_reg_3144_pp0_iter71_reg <= p_read_40_reg_3144_pp0_iter70_reg;
            p_read_40_reg_3144_pp0_iter72_reg <= p_read_40_reg_3144_pp0_iter71_reg;
            p_read_40_reg_3144_pp0_iter73_reg <= p_read_40_reg_3144_pp0_iter72_reg;
            p_read_40_reg_3144_pp0_iter74_reg <= p_read_40_reg_3144_pp0_iter73_reg;
            p_read_40_reg_3144_pp0_iter75_reg <= p_read_40_reg_3144_pp0_iter74_reg;
            p_read_40_reg_3144_pp0_iter76_reg <= p_read_40_reg_3144_pp0_iter75_reg;
            p_read_40_reg_3144_pp0_iter7_reg <= p_read_40_reg_3144_pp0_iter6_reg;
            p_read_40_reg_3144_pp0_iter8_reg <= p_read_40_reg_3144_pp0_iter7_reg;
            p_read_40_reg_3144_pp0_iter9_reg <= p_read_40_reg_3144_pp0_iter8_reg;
            p_read_41_reg_3149 <= p_read23_int_reg;
            p_read_41_reg_3149_pp0_iter10_reg <= p_read_41_reg_3149_pp0_iter9_reg;
            p_read_41_reg_3149_pp0_iter11_reg <= p_read_41_reg_3149_pp0_iter10_reg;
            p_read_41_reg_3149_pp0_iter12_reg <= p_read_41_reg_3149_pp0_iter11_reg;
            p_read_41_reg_3149_pp0_iter13_reg <= p_read_41_reg_3149_pp0_iter12_reg;
            p_read_41_reg_3149_pp0_iter14_reg <= p_read_41_reg_3149_pp0_iter13_reg;
            p_read_41_reg_3149_pp0_iter15_reg <= p_read_41_reg_3149_pp0_iter14_reg;
            p_read_41_reg_3149_pp0_iter16_reg <= p_read_41_reg_3149_pp0_iter15_reg;
            p_read_41_reg_3149_pp0_iter17_reg <= p_read_41_reg_3149_pp0_iter16_reg;
            p_read_41_reg_3149_pp0_iter18_reg <= p_read_41_reg_3149_pp0_iter17_reg;
            p_read_41_reg_3149_pp0_iter19_reg <= p_read_41_reg_3149_pp0_iter18_reg;
            p_read_41_reg_3149_pp0_iter1_reg <= p_read_41_reg_3149;
            p_read_41_reg_3149_pp0_iter20_reg <= p_read_41_reg_3149_pp0_iter19_reg;
            p_read_41_reg_3149_pp0_iter21_reg <= p_read_41_reg_3149_pp0_iter20_reg;
            p_read_41_reg_3149_pp0_iter22_reg <= p_read_41_reg_3149_pp0_iter21_reg;
            p_read_41_reg_3149_pp0_iter23_reg <= p_read_41_reg_3149_pp0_iter22_reg;
            p_read_41_reg_3149_pp0_iter24_reg <= p_read_41_reg_3149_pp0_iter23_reg;
            p_read_41_reg_3149_pp0_iter25_reg <= p_read_41_reg_3149_pp0_iter24_reg;
            p_read_41_reg_3149_pp0_iter26_reg <= p_read_41_reg_3149_pp0_iter25_reg;
            p_read_41_reg_3149_pp0_iter27_reg <= p_read_41_reg_3149_pp0_iter26_reg;
            p_read_41_reg_3149_pp0_iter28_reg <= p_read_41_reg_3149_pp0_iter27_reg;
            p_read_41_reg_3149_pp0_iter29_reg <= p_read_41_reg_3149_pp0_iter28_reg;
            p_read_41_reg_3149_pp0_iter2_reg <= p_read_41_reg_3149_pp0_iter1_reg;
            p_read_41_reg_3149_pp0_iter30_reg <= p_read_41_reg_3149_pp0_iter29_reg;
            p_read_41_reg_3149_pp0_iter31_reg <= p_read_41_reg_3149_pp0_iter30_reg;
            p_read_41_reg_3149_pp0_iter32_reg <= p_read_41_reg_3149_pp0_iter31_reg;
            p_read_41_reg_3149_pp0_iter33_reg <= p_read_41_reg_3149_pp0_iter32_reg;
            p_read_41_reg_3149_pp0_iter34_reg <= p_read_41_reg_3149_pp0_iter33_reg;
            p_read_41_reg_3149_pp0_iter35_reg <= p_read_41_reg_3149_pp0_iter34_reg;
            p_read_41_reg_3149_pp0_iter36_reg <= p_read_41_reg_3149_pp0_iter35_reg;
            p_read_41_reg_3149_pp0_iter37_reg <= p_read_41_reg_3149_pp0_iter36_reg;
            p_read_41_reg_3149_pp0_iter38_reg <= p_read_41_reg_3149_pp0_iter37_reg;
            p_read_41_reg_3149_pp0_iter39_reg <= p_read_41_reg_3149_pp0_iter38_reg;
            p_read_41_reg_3149_pp0_iter3_reg <= p_read_41_reg_3149_pp0_iter2_reg;
            p_read_41_reg_3149_pp0_iter40_reg <= p_read_41_reg_3149_pp0_iter39_reg;
            p_read_41_reg_3149_pp0_iter41_reg <= p_read_41_reg_3149_pp0_iter40_reg;
            p_read_41_reg_3149_pp0_iter42_reg <= p_read_41_reg_3149_pp0_iter41_reg;
            p_read_41_reg_3149_pp0_iter43_reg <= p_read_41_reg_3149_pp0_iter42_reg;
            p_read_41_reg_3149_pp0_iter44_reg <= p_read_41_reg_3149_pp0_iter43_reg;
            p_read_41_reg_3149_pp0_iter45_reg <= p_read_41_reg_3149_pp0_iter44_reg;
            p_read_41_reg_3149_pp0_iter46_reg <= p_read_41_reg_3149_pp0_iter45_reg;
            p_read_41_reg_3149_pp0_iter47_reg <= p_read_41_reg_3149_pp0_iter46_reg;
            p_read_41_reg_3149_pp0_iter48_reg <= p_read_41_reg_3149_pp0_iter47_reg;
            p_read_41_reg_3149_pp0_iter49_reg <= p_read_41_reg_3149_pp0_iter48_reg;
            p_read_41_reg_3149_pp0_iter4_reg <= p_read_41_reg_3149_pp0_iter3_reg;
            p_read_41_reg_3149_pp0_iter50_reg <= p_read_41_reg_3149_pp0_iter49_reg;
            p_read_41_reg_3149_pp0_iter51_reg <= p_read_41_reg_3149_pp0_iter50_reg;
            p_read_41_reg_3149_pp0_iter52_reg <= p_read_41_reg_3149_pp0_iter51_reg;
            p_read_41_reg_3149_pp0_iter53_reg <= p_read_41_reg_3149_pp0_iter52_reg;
            p_read_41_reg_3149_pp0_iter54_reg <= p_read_41_reg_3149_pp0_iter53_reg;
            p_read_41_reg_3149_pp0_iter55_reg <= p_read_41_reg_3149_pp0_iter54_reg;
            p_read_41_reg_3149_pp0_iter56_reg <= p_read_41_reg_3149_pp0_iter55_reg;
            p_read_41_reg_3149_pp0_iter57_reg <= p_read_41_reg_3149_pp0_iter56_reg;
            p_read_41_reg_3149_pp0_iter58_reg <= p_read_41_reg_3149_pp0_iter57_reg;
            p_read_41_reg_3149_pp0_iter59_reg <= p_read_41_reg_3149_pp0_iter58_reg;
            p_read_41_reg_3149_pp0_iter5_reg <= p_read_41_reg_3149_pp0_iter4_reg;
            p_read_41_reg_3149_pp0_iter60_reg <= p_read_41_reg_3149_pp0_iter59_reg;
            p_read_41_reg_3149_pp0_iter61_reg <= p_read_41_reg_3149_pp0_iter60_reg;
            p_read_41_reg_3149_pp0_iter62_reg <= p_read_41_reg_3149_pp0_iter61_reg;
            p_read_41_reg_3149_pp0_iter63_reg <= p_read_41_reg_3149_pp0_iter62_reg;
            p_read_41_reg_3149_pp0_iter64_reg <= p_read_41_reg_3149_pp0_iter63_reg;
            p_read_41_reg_3149_pp0_iter65_reg <= p_read_41_reg_3149_pp0_iter64_reg;
            p_read_41_reg_3149_pp0_iter66_reg <= p_read_41_reg_3149_pp0_iter65_reg;
            p_read_41_reg_3149_pp0_iter67_reg <= p_read_41_reg_3149_pp0_iter66_reg;
            p_read_41_reg_3149_pp0_iter68_reg <= p_read_41_reg_3149_pp0_iter67_reg;
            p_read_41_reg_3149_pp0_iter69_reg <= p_read_41_reg_3149_pp0_iter68_reg;
            p_read_41_reg_3149_pp0_iter6_reg <= p_read_41_reg_3149_pp0_iter5_reg;
            p_read_41_reg_3149_pp0_iter70_reg <= p_read_41_reg_3149_pp0_iter69_reg;
            p_read_41_reg_3149_pp0_iter71_reg <= p_read_41_reg_3149_pp0_iter70_reg;
            p_read_41_reg_3149_pp0_iter72_reg <= p_read_41_reg_3149_pp0_iter71_reg;
            p_read_41_reg_3149_pp0_iter73_reg <= p_read_41_reg_3149_pp0_iter72_reg;
            p_read_41_reg_3149_pp0_iter74_reg <= p_read_41_reg_3149_pp0_iter73_reg;
            p_read_41_reg_3149_pp0_iter75_reg <= p_read_41_reg_3149_pp0_iter74_reg;
            p_read_41_reg_3149_pp0_iter76_reg <= p_read_41_reg_3149_pp0_iter75_reg;
            p_read_41_reg_3149_pp0_iter7_reg <= p_read_41_reg_3149_pp0_iter6_reg;
            p_read_41_reg_3149_pp0_iter8_reg <= p_read_41_reg_3149_pp0_iter7_reg;
            p_read_41_reg_3149_pp0_iter9_reg <= p_read_41_reg_3149_pp0_iter8_reg;
            p_read_42_reg_3154 <= p_read22_int_reg;
            p_read_42_reg_3154_pp0_iter10_reg <= p_read_42_reg_3154_pp0_iter9_reg;
            p_read_42_reg_3154_pp0_iter11_reg <= p_read_42_reg_3154_pp0_iter10_reg;
            p_read_42_reg_3154_pp0_iter12_reg <= p_read_42_reg_3154_pp0_iter11_reg;
            p_read_42_reg_3154_pp0_iter13_reg <= p_read_42_reg_3154_pp0_iter12_reg;
            p_read_42_reg_3154_pp0_iter14_reg <= p_read_42_reg_3154_pp0_iter13_reg;
            p_read_42_reg_3154_pp0_iter15_reg <= p_read_42_reg_3154_pp0_iter14_reg;
            p_read_42_reg_3154_pp0_iter16_reg <= p_read_42_reg_3154_pp0_iter15_reg;
            p_read_42_reg_3154_pp0_iter17_reg <= p_read_42_reg_3154_pp0_iter16_reg;
            p_read_42_reg_3154_pp0_iter18_reg <= p_read_42_reg_3154_pp0_iter17_reg;
            p_read_42_reg_3154_pp0_iter19_reg <= p_read_42_reg_3154_pp0_iter18_reg;
            p_read_42_reg_3154_pp0_iter1_reg <= p_read_42_reg_3154;
            p_read_42_reg_3154_pp0_iter20_reg <= p_read_42_reg_3154_pp0_iter19_reg;
            p_read_42_reg_3154_pp0_iter21_reg <= p_read_42_reg_3154_pp0_iter20_reg;
            p_read_42_reg_3154_pp0_iter22_reg <= p_read_42_reg_3154_pp0_iter21_reg;
            p_read_42_reg_3154_pp0_iter23_reg <= p_read_42_reg_3154_pp0_iter22_reg;
            p_read_42_reg_3154_pp0_iter24_reg <= p_read_42_reg_3154_pp0_iter23_reg;
            p_read_42_reg_3154_pp0_iter25_reg <= p_read_42_reg_3154_pp0_iter24_reg;
            p_read_42_reg_3154_pp0_iter26_reg <= p_read_42_reg_3154_pp0_iter25_reg;
            p_read_42_reg_3154_pp0_iter27_reg <= p_read_42_reg_3154_pp0_iter26_reg;
            p_read_42_reg_3154_pp0_iter28_reg <= p_read_42_reg_3154_pp0_iter27_reg;
            p_read_42_reg_3154_pp0_iter29_reg <= p_read_42_reg_3154_pp0_iter28_reg;
            p_read_42_reg_3154_pp0_iter2_reg <= p_read_42_reg_3154_pp0_iter1_reg;
            p_read_42_reg_3154_pp0_iter30_reg <= p_read_42_reg_3154_pp0_iter29_reg;
            p_read_42_reg_3154_pp0_iter31_reg <= p_read_42_reg_3154_pp0_iter30_reg;
            p_read_42_reg_3154_pp0_iter32_reg <= p_read_42_reg_3154_pp0_iter31_reg;
            p_read_42_reg_3154_pp0_iter33_reg <= p_read_42_reg_3154_pp0_iter32_reg;
            p_read_42_reg_3154_pp0_iter34_reg <= p_read_42_reg_3154_pp0_iter33_reg;
            p_read_42_reg_3154_pp0_iter35_reg <= p_read_42_reg_3154_pp0_iter34_reg;
            p_read_42_reg_3154_pp0_iter36_reg <= p_read_42_reg_3154_pp0_iter35_reg;
            p_read_42_reg_3154_pp0_iter37_reg <= p_read_42_reg_3154_pp0_iter36_reg;
            p_read_42_reg_3154_pp0_iter38_reg <= p_read_42_reg_3154_pp0_iter37_reg;
            p_read_42_reg_3154_pp0_iter39_reg <= p_read_42_reg_3154_pp0_iter38_reg;
            p_read_42_reg_3154_pp0_iter3_reg <= p_read_42_reg_3154_pp0_iter2_reg;
            p_read_42_reg_3154_pp0_iter40_reg <= p_read_42_reg_3154_pp0_iter39_reg;
            p_read_42_reg_3154_pp0_iter41_reg <= p_read_42_reg_3154_pp0_iter40_reg;
            p_read_42_reg_3154_pp0_iter42_reg <= p_read_42_reg_3154_pp0_iter41_reg;
            p_read_42_reg_3154_pp0_iter43_reg <= p_read_42_reg_3154_pp0_iter42_reg;
            p_read_42_reg_3154_pp0_iter44_reg <= p_read_42_reg_3154_pp0_iter43_reg;
            p_read_42_reg_3154_pp0_iter45_reg <= p_read_42_reg_3154_pp0_iter44_reg;
            p_read_42_reg_3154_pp0_iter46_reg <= p_read_42_reg_3154_pp0_iter45_reg;
            p_read_42_reg_3154_pp0_iter47_reg <= p_read_42_reg_3154_pp0_iter46_reg;
            p_read_42_reg_3154_pp0_iter48_reg <= p_read_42_reg_3154_pp0_iter47_reg;
            p_read_42_reg_3154_pp0_iter49_reg <= p_read_42_reg_3154_pp0_iter48_reg;
            p_read_42_reg_3154_pp0_iter4_reg <= p_read_42_reg_3154_pp0_iter3_reg;
            p_read_42_reg_3154_pp0_iter50_reg <= p_read_42_reg_3154_pp0_iter49_reg;
            p_read_42_reg_3154_pp0_iter51_reg <= p_read_42_reg_3154_pp0_iter50_reg;
            p_read_42_reg_3154_pp0_iter52_reg <= p_read_42_reg_3154_pp0_iter51_reg;
            p_read_42_reg_3154_pp0_iter53_reg <= p_read_42_reg_3154_pp0_iter52_reg;
            p_read_42_reg_3154_pp0_iter54_reg <= p_read_42_reg_3154_pp0_iter53_reg;
            p_read_42_reg_3154_pp0_iter55_reg <= p_read_42_reg_3154_pp0_iter54_reg;
            p_read_42_reg_3154_pp0_iter56_reg <= p_read_42_reg_3154_pp0_iter55_reg;
            p_read_42_reg_3154_pp0_iter57_reg <= p_read_42_reg_3154_pp0_iter56_reg;
            p_read_42_reg_3154_pp0_iter58_reg <= p_read_42_reg_3154_pp0_iter57_reg;
            p_read_42_reg_3154_pp0_iter59_reg <= p_read_42_reg_3154_pp0_iter58_reg;
            p_read_42_reg_3154_pp0_iter5_reg <= p_read_42_reg_3154_pp0_iter4_reg;
            p_read_42_reg_3154_pp0_iter60_reg <= p_read_42_reg_3154_pp0_iter59_reg;
            p_read_42_reg_3154_pp0_iter61_reg <= p_read_42_reg_3154_pp0_iter60_reg;
            p_read_42_reg_3154_pp0_iter62_reg <= p_read_42_reg_3154_pp0_iter61_reg;
            p_read_42_reg_3154_pp0_iter63_reg <= p_read_42_reg_3154_pp0_iter62_reg;
            p_read_42_reg_3154_pp0_iter64_reg <= p_read_42_reg_3154_pp0_iter63_reg;
            p_read_42_reg_3154_pp0_iter65_reg <= p_read_42_reg_3154_pp0_iter64_reg;
            p_read_42_reg_3154_pp0_iter66_reg <= p_read_42_reg_3154_pp0_iter65_reg;
            p_read_42_reg_3154_pp0_iter67_reg <= p_read_42_reg_3154_pp0_iter66_reg;
            p_read_42_reg_3154_pp0_iter68_reg <= p_read_42_reg_3154_pp0_iter67_reg;
            p_read_42_reg_3154_pp0_iter69_reg <= p_read_42_reg_3154_pp0_iter68_reg;
            p_read_42_reg_3154_pp0_iter6_reg <= p_read_42_reg_3154_pp0_iter5_reg;
            p_read_42_reg_3154_pp0_iter70_reg <= p_read_42_reg_3154_pp0_iter69_reg;
            p_read_42_reg_3154_pp0_iter71_reg <= p_read_42_reg_3154_pp0_iter70_reg;
            p_read_42_reg_3154_pp0_iter72_reg <= p_read_42_reg_3154_pp0_iter71_reg;
            p_read_42_reg_3154_pp0_iter73_reg <= p_read_42_reg_3154_pp0_iter72_reg;
            p_read_42_reg_3154_pp0_iter74_reg <= p_read_42_reg_3154_pp0_iter73_reg;
            p_read_42_reg_3154_pp0_iter75_reg <= p_read_42_reg_3154_pp0_iter74_reg;
            p_read_42_reg_3154_pp0_iter76_reg <= p_read_42_reg_3154_pp0_iter75_reg;
            p_read_42_reg_3154_pp0_iter7_reg <= p_read_42_reg_3154_pp0_iter6_reg;
            p_read_42_reg_3154_pp0_iter8_reg <= p_read_42_reg_3154_pp0_iter7_reg;
            p_read_42_reg_3154_pp0_iter9_reg <= p_read_42_reg_3154_pp0_iter8_reg;
            p_read_43_reg_3159 <= p_read21_int_reg;
            p_read_43_reg_3159_pp0_iter10_reg <= p_read_43_reg_3159_pp0_iter9_reg;
            p_read_43_reg_3159_pp0_iter11_reg <= p_read_43_reg_3159_pp0_iter10_reg;
            p_read_43_reg_3159_pp0_iter12_reg <= p_read_43_reg_3159_pp0_iter11_reg;
            p_read_43_reg_3159_pp0_iter13_reg <= p_read_43_reg_3159_pp0_iter12_reg;
            p_read_43_reg_3159_pp0_iter14_reg <= p_read_43_reg_3159_pp0_iter13_reg;
            p_read_43_reg_3159_pp0_iter15_reg <= p_read_43_reg_3159_pp0_iter14_reg;
            p_read_43_reg_3159_pp0_iter16_reg <= p_read_43_reg_3159_pp0_iter15_reg;
            p_read_43_reg_3159_pp0_iter17_reg <= p_read_43_reg_3159_pp0_iter16_reg;
            p_read_43_reg_3159_pp0_iter18_reg <= p_read_43_reg_3159_pp0_iter17_reg;
            p_read_43_reg_3159_pp0_iter19_reg <= p_read_43_reg_3159_pp0_iter18_reg;
            p_read_43_reg_3159_pp0_iter1_reg <= p_read_43_reg_3159;
            p_read_43_reg_3159_pp0_iter20_reg <= p_read_43_reg_3159_pp0_iter19_reg;
            p_read_43_reg_3159_pp0_iter21_reg <= p_read_43_reg_3159_pp0_iter20_reg;
            p_read_43_reg_3159_pp0_iter22_reg <= p_read_43_reg_3159_pp0_iter21_reg;
            p_read_43_reg_3159_pp0_iter23_reg <= p_read_43_reg_3159_pp0_iter22_reg;
            p_read_43_reg_3159_pp0_iter24_reg <= p_read_43_reg_3159_pp0_iter23_reg;
            p_read_43_reg_3159_pp0_iter25_reg <= p_read_43_reg_3159_pp0_iter24_reg;
            p_read_43_reg_3159_pp0_iter26_reg <= p_read_43_reg_3159_pp0_iter25_reg;
            p_read_43_reg_3159_pp0_iter27_reg <= p_read_43_reg_3159_pp0_iter26_reg;
            p_read_43_reg_3159_pp0_iter28_reg <= p_read_43_reg_3159_pp0_iter27_reg;
            p_read_43_reg_3159_pp0_iter29_reg <= p_read_43_reg_3159_pp0_iter28_reg;
            p_read_43_reg_3159_pp0_iter2_reg <= p_read_43_reg_3159_pp0_iter1_reg;
            p_read_43_reg_3159_pp0_iter30_reg <= p_read_43_reg_3159_pp0_iter29_reg;
            p_read_43_reg_3159_pp0_iter31_reg <= p_read_43_reg_3159_pp0_iter30_reg;
            p_read_43_reg_3159_pp0_iter32_reg <= p_read_43_reg_3159_pp0_iter31_reg;
            p_read_43_reg_3159_pp0_iter33_reg <= p_read_43_reg_3159_pp0_iter32_reg;
            p_read_43_reg_3159_pp0_iter34_reg <= p_read_43_reg_3159_pp0_iter33_reg;
            p_read_43_reg_3159_pp0_iter35_reg <= p_read_43_reg_3159_pp0_iter34_reg;
            p_read_43_reg_3159_pp0_iter36_reg <= p_read_43_reg_3159_pp0_iter35_reg;
            p_read_43_reg_3159_pp0_iter37_reg <= p_read_43_reg_3159_pp0_iter36_reg;
            p_read_43_reg_3159_pp0_iter38_reg <= p_read_43_reg_3159_pp0_iter37_reg;
            p_read_43_reg_3159_pp0_iter39_reg <= p_read_43_reg_3159_pp0_iter38_reg;
            p_read_43_reg_3159_pp0_iter3_reg <= p_read_43_reg_3159_pp0_iter2_reg;
            p_read_43_reg_3159_pp0_iter40_reg <= p_read_43_reg_3159_pp0_iter39_reg;
            p_read_43_reg_3159_pp0_iter41_reg <= p_read_43_reg_3159_pp0_iter40_reg;
            p_read_43_reg_3159_pp0_iter42_reg <= p_read_43_reg_3159_pp0_iter41_reg;
            p_read_43_reg_3159_pp0_iter43_reg <= p_read_43_reg_3159_pp0_iter42_reg;
            p_read_43_reg_3159_pp0_iter44_reg <= p_read_43_reg_3159_pp0_iter43_reg;
            p_read_43_reg_3159_pp0_iter45_reg <= p_read_43_reg_3159_pp0_iter44_reg;
            p_read_43_reg_3159_pp0_iter46_reg <= p_read_43_reg_3159_pp0_iter45_reg;
            p_read_43_reg_3159_pp0_iter47_reg <= p_read_43_reg_3159_pp0_iter46_reg;
            p_read_43_reg_3159_pp0_iter48_reg <= p_read_43_reg_3159_pp0_iter47_reg;
            p_read_43_reg_3159_pp0_iter49_reg <= p_read_43_reg_3159_pp0_iter48_reg;
            p_read_43_reg_3159_pp0_iter4_reg <= p_read_43_reg_3159_pp0_iter3_reg;
            p_read_43_reg_3159_pp0_iter50_reg <= p_read_43_reg_3159_pp0_iter49_reg;
            p_read_43_reg_3159_pp0_iter51_reg <= p_read_43_reg_3159_pp0_iter50_reg;
            p_read_43_reg_3159_pp0_iter52_reg <= p_read_43_reg_3159_pp0_iter51_reg;
            p_read_43_reg_3159_pp0_iter53_reg <= p_read_43_reg_3159_pp0_iter52_reg;
            p_read_43_reg_3159_pp0_iter54_reg <= p_read_43_reg_3159_pp0_iter53_reg;
            p_read_43_reg_3159_pp0_iter55_reg <= p_read_43_reg_3159_pp0_iter54_reg;
            p_read_43_reg_3159_pp0_iter56_reg <= p_read_43_reg_3159_pp0_iter55_reg;
            p_read_43_reg_3159_pp0_iter57_reg <= p_read_43_reg_3159_pp0_iter56_reg;
            p_read_43_reg_3159_pp0_iter58_reg <= p_read_43_reg_3159_pp0_iter57_reg;
            p_read_43_reg_3159_pp0_iter59_reg <= p_read_43_reg_3159_pp0_iter58_reg;
            p_read_43_reg_3159_pp0_iter5_reg <= p_read_43_reg_3159_pp0_iter4_reg;
            p_read_43_reg_3159_pp0_iter60_reg <= p_read_43_reg_3159_pp0_iter59_reg;
            p_read_43_reg_3159_pp0_iter61_reg <= p_read_43_reg_3159_pp0_iter60_reg;
            p_read_43_reg_3159_pp0_iter62_reg <= p_read_43_reg_3159_pp0_iter61_reg;
            p_read_43_reg_3159_pp0_iter63_reg <= p_read_43_reg_3159_pp0_iter62_reg;
            p_read_43_reg_3159_pp0_iter64_reg <= p_read_43_reg_3159_pp0_iter63_reg;
            p_read_43_reg_3159_pp0_iter65_reg <= p_read_43_reg_3159_pp0_iter64_reg;
            p_read_43_reg_3159_pp0_iter66_reg <= p_read_43_reg_3159_pp0_iter65_reg;
            p_read_43_reg_3159_pp0_iter67_reg <= p_read_43_reg_3159_pp0_iter66_reg;
            p_read_43_reg_3159_pp0_iter68_reg <= p_read_43_reg_3159_pp0_iter67_reg;
            p_read_43_reg_3159_pp0_iter69_reg <= p_read_43_reg_3159_pp0_iter68_reg;
            p_read_43_reg_3159_pp0_iter6_reg <= p_read_43_reg_3159_pp0_iter5_reg;
            p_read_43_reg_3159_pp0_iter70_reg <= p_read_43_reg_3159_pp0_iter69_reg;
            p_read_43_reg_3159_pp0_iter71_reg <= p_read_43_reg_3159_pp0_iter70_reg;
            p_read_43_reg_3159_pp0_iter72_reg <= p_read_43_reg_3159_pp0_iter71_reg;
            p_read_43_reg_3159_pp0_iter73_reg <= p_read_43_reg_3159_pp0_iter72_reg;
            p_read_43_reg_3159_pp0_iter74_reg <= p_read_43_reg_3159_pp0_iter73_reg;
            p_read_43_reg_3159_pp0_iter75_reg <= p_read_43_reg_3159_pp0_iter74_reg;
            p_read_43_reg_3159_pp0_iter76_reg <= p_read_43_reg_3159_pp0_iter75_reg;
            p_read_43_reg_3159_pp0_iter7_reg <= p_read_43_reg_3159_pp0_iter6_reg;
            p_read_43_reg_3159_pp0_iter8_reg <= p_read_43_reg_3159_pp0_iter7_reg;
            p_read_43_reg_3159_pp0_iter9_reg <= p_read_43_reg_3159_pp0_iter8_reg;
            p_read_44_reg_3164 <= p_read20_int_reg;
            p_read_44_reg_3164_pp0_iter10_reg <= p_read_44_reg_3164_pp0_iter9_reg;
            p_read_44_reg_3164_pp0_iter11_reg <= p_read_44_reg_3164_pp0_iter10_reg;
            p_read_44_reg_3164_pp0_iter12_reg <= p_read_44_reg_3164_pp0_iter11_reg;
            p_read_44_reg_3164_pp0_iter13_reg <= p_read_44_reg_3164_pp0_iter12_reg;
            p_read_44_reg_3164_pp0_iter14_reg <= p_read_44_reg_3164_pp0_iter13_reg;
            p_read_44_reg_3164_pp0_iter15_reg <= p_read_44_reg_3164_pp0_iter14_reg;
            p_read_44_reg_3164_pp0_iter16_reg <= p_read_44_reg_3164_pp0_iter15_reg;
            p_read_44_reg_3164_pp0_iter17_reg <= p_read_44_reg_3164_pp0_iter16_reg;
            p_read_44_reg_3164_pp0_iter18_reg <= p_read_44_reg_3164_pp0_iter17_reg;
            p_read_44_reg_3164_pp0_iter19_reg <= p_read_44_reg_3164_pp0_iter18_reg;
            p_read_44_reg_3164_pp0_iter1_reg <= p_read_44_reg_3164;
            p_read_44_reg_3164_pp0_iter20_reg <= p_read_44_reg_3164_pp0_iter19_reg;
            p_read_44_reg_3164_pp0_iter21_reg <= p_read_44_reg_3164_pp0_iter20_reg;
            p_read_44_reg_3164_pp0_iter22_reg <= p_read_44_reg_3164_pp0_iter21_reg;
            p_read_44_reg_3164_pp0_iter23_reg <= p_read_44_reg_3164_pp0_iter22_reg;
            p_read_44_reg_3164_pp0_iter24_reg <= p_read_44_reg_3164_pp0_iter23_reg;
            p_read_44_reg_3164_pp0_iter25_reg <= p_read_44_reg_3164_pp0_iter24_reg;
            p_read_44_reg_3164_pp0_iter26_reg <= p_read_44_reg_3164_pp0_iter25_reg;
            p_read_44_reg_3164_pp0_iter27_reg <= p_read_44_reg_3164_pp0_iter26_reg;
            p_read_44_reg_3164_pp0_iter28_reg <= p_read_44_reg_3164_pp0_iter27_reg;
            p_read_44_reg_3164_pp0_iter29_reg <= p_read_44_reg_3164_pp0_iter28_reg;
            p_read_44_reg_3164_pp0_iter2_reg <= p_read_44_reg_3164_pp0_iter1_reg;
            p_read_44_reg_3164_pp0_iter30_reg <= p_read_44_reg_3164_pp0_iter29_reg;
            p_read_44_reg_3164_pp0_iter31_reg <= p_read_44_reg_3164_pp0_iter30_reg;
            p_read_44_reg_3164_pp0_iter32_reg <= p_read_44_reg_3164_pp0_iter31_reg;
            p_read_44_reg_3164_pp0_iter33_reg <= p_read_44_reg_3164_pp0_iter32_reg;
            p_read_44_reg_3164_pp0_iter34_reg <= p_read_44_reg_3164_pp0_iter33_reg;
            p_read_44_reg_3164_pp0_iter35_reg <= p_read_44_reg_3164_pp0_iter34_reg;
            p_read_44_reg_3164_pp0_iter36_reg <= p_read_44_reg_3164_pp0_iter35_reg;
            p_read_44_reg_3164_pp0_iter37_reg <= p_read_44_reg_3164_pp0_iter36_reg;
            p_read_44_reg_3164_pp0_iter38_reg <= p_read_44_reg_3164_pp0_iter37_reg;
            p_read_44_reg_3164_pp0_iter39_reg <= p_read_44_reg_3164_pp0_iter38_reg;
            p_read_44_reg_3164_pp0_iter3_reg <= p_read_44_reg_3164_pp0_iter2_reg;
            p_read_44_reg_3164_pp0_iter40_reg <= p_read_44_reg_3164_pp0_iter39_reg;
            p_read_44_reg_3164_pp0_iter41_reg <= p_read_44_reg_3164_pp0_iter40_reg;
            p_read_44_reg_3164_pp0_iter42_reg <= p_read_44_reg_3164_pp0_iter41_reg;
            p_read_44_reg_3164_pp0_iter43_reg <= p_read_44_reg_3164_pp0_iter42_reg;
            p_read_44_reg_3164_pp0_iter44_reg <= p_read_44_reg_3164_pp0_iter43_reg;
            p_read_44_reg_3164_pp0_iter45_reg <= p_read_44_reg_3164_pp0_iter44_reg;
            p_read_44_reg_3164_pp0_iter46_reg <= p_read_44_reg_3164_pp0_iter45_reg;
            p_read_44_reg_3164_pp0_iter47_reg <= p_read_44_reg_3164_pp0_iter46_reg;
            p_read_44_reg_3164_pp0_iter48_reg <= p_read_44_reg_3164_pp0_iter47_reg;
            p_read_44_reg_3164_pp0_iter49_reg <= p_read_44_reg_3164_pp0_iter48_reg;
            p_read_44_reg_3164_pp0_iter4_reg <= p_read_44_reg_3164_pp0_iter3_reg;
            p_read_44_reg_3164_pp0_iter50_reg <= p_read_44_reg_3164_pp0_iter49_reg;
            p_read_44_reg_3164_pp0_iter51_reg <= p_read_44_reg_3164_pp0_iter50_reg;
            p_read_44_reg_3164_pp0_iter52_reg <= p_read_44_reg_3164_pp0_iter51_reg;
            p_read_44_reg_3164_pp0_iter53_reg <= p_read_44_reg_3164_pp0_iter52_reg;
            p_read_44_reg_3164_pp0_iter54_reg <= p_read_44_reg_3164_pp0_iter53_reg;
            p_read_44_reg_3164_pp0_iter55_reg <= p_read_44_reg_3164_pp0_iter54_reg;
            p_read_44_reg_3164_pp0_iter56_reg <= p_read_44_reg_3164_pp0_iter55_reg;
            p_read_44_reg_3164_pp0_iter57_reg <= p_read_44_reg_3164_pp0_iter56_reg;
            p_read_44_reg_3164_pp0_iter58_reg <= p_read_44_reg_3164_pp0_iter57_reg;
            p_read_44_reg_3164_pp0_iter59_reg <= p_read_44_reg_3164_pp0_iter58_reg;
            p_read_44_reg_3164_pp0_iter5_reg <= p_read_44_reg_3164_pp0_iter4_reg;
            p_read_44_reg_3164_pp0_iter60_reg <= p_read_44_reg_3164_pp0_iter59_reg;
            p_read_44_reg_3164_pp0_iter61_reg <= p_read_44_reg_3164_pp0_iter60_reg;
            p_read_44_reg_3164_pp0_iter62_reg <= p_read_44_reg_3164_pp0_iter61_reg;
            p_read_44_reg_3164_pp0_iter63_reg <= p_read_44_reg_3164_pp0_iter62_reg;
            p_read_44_reg_3164_pp0_iter64_reg <= p_read_44_reg_3164_pp0_iter63_reg;
            p_read_44_reg_3164_pp0_iter65_reg <= p_read_44_reg_3164_pp0_iter64_reg;
            p_read_44_reg_3164_pp0_iter66_reg <= p_read_44_reg_3164_pp0_iter65_reg;
            p_read_44_reg_3164_pp0_iter67_reg <= p_read_44_reg_3164_pp0_iter66_reg;
            p_read_44_reg_3164_pp0_iter68_reg <= p_read_44_reg_3164_pp0_iter67_reg;
            p_read_44_reg_3164_pp0_iter69_reg <= p_read_44_reg_3164_pp0_iter68_reg;
            p_read_44_reg_3164_pp0_iter6_reg <= p_read_44_reg_3164_pp0_iter5_reg;
            p_read_44_reg_3164_pp0_iter70_reg <= p_read_44_reg_3164_pp0_iter69_reg;
            p_read_44_reg_3164_pp0_iter71_reg <= p_read_44_reg_3164_pp0_iter70_reg;
            p_read_44_reg_3164_pp0_iter72_reg <= p_read_44_reg_3164_pp0_iter71_reg;
            p_read_44_reg_3164_pp0_iter73_reg <= p_read_44_reg_3164_pp0_iter72_reg;
            p_read_44_reg_3164_pp0_iter74_reg <= p_read_44_reg_3164_pp0_iter73_reg;
            p_read_44_reg_3164_pp0_iter75_reg <= p_read_44_reg_3164_pp0_iter74_reg;
            p_read_44_reg_3164_pp0_iter76_reg <= p_read_44_reg_3164_pp0_iter75_reg;
            p_read_44_reg_3164_pp0_iter7_reg <= p_read_44_reg_3164_pp0_iter6_reg;
            p_read_44_reg_3164_pp0_iter8_reg <= p_read_44_reg_3164_pp0_iter7_reg;
            p_read_44_reg_3164_pp0_iter9_reg <= p_read_44_reg_3164_pp0_iter8_reg;
            p_read_45_reg_3169 <= p_read19_int_reg;
            p_read_45_reg_3169_pp0_iter10_reg <= p_read_45_reg_3169_pp0_iter9_reg;
            p_read_45_reg_3169_pp0_iter11_reg <= p_read_45_reg_3169_pp0_iter10_reg;
            p_read_45_reg_3169_pp0_iter12_reg <= p_read_45_reg_3169_pp0_iter11_reg;
            p_read_45_reg_3169_pp0_iter13_reg <= p_read_45_reg_3169_pp0_iter12_reg;
            p_read_45_reg_3169_pp0_iter14_reg <= p_read_45_reg_3169_pp0_iter13_reg;
            p_read_45_reg_3169_pp0_iter15_reg <= p_read_45_reg_3169_pp0_iter14_reg;
            p_read_45_reg_3169_pp0_iter16_reg <= p_read_45_reg_3169_pp0_iter15_reg;
            p_read_45_reg_3169_pp0_iter17_reg <= p_read_45_reg_3169_pp0_iter16_reg;
            p_read_45_reg_3169_pp0_iter18_reg <= p_read_45_reg_3169_pp0_iter17_reg;
            p_read_45_reg_3169_pp0_iter19_reg <= p_read_45_reg_3169_pp0_iter18_reg;
            p_read_45_reg_3169_pp0_iter1_reg <= p_read_45_reg_3169;
            p_read_45_reg_3169_pp0_iter20_reg <= p_read_45_reg_3169_pp0_iter19_reg;
            p_read_45_reg_3169_pp0_iter21_reg <= p_read_45_reg_3169_pp0_iter20_reg;
            p_read_45_reg_3169_pp0_iter22_reg <= p_read_45_reg_3169_pp0_iter21_reg;
            p_read_45_reg_3169_pp0_iter23_reg <= p_read_45_reg_3169_pp0_iter22_reg;
            p_read_45_reg_3169_pp0_iter24_reg <= p_read_45_reg_3169_pp0_iter23_reg;
            p_read_45_reg_3169_pp0_iter25_reg <= p_read_45_reg_3169_pp0_iter24_reg;
            p_read_45_reg_3169_pp0_iter26_reg <= p_read_45_reg_3169_pp0_iter25_reg;
            p_read_45_reg_3169_pp0_iter27_reg <= p_read_45_reg_3169_pp0_iter26_reg;
            p_read_45_reg_3169_pp0_iter28_reg <= p_read_45_reg_3169_pp0_iter27_reg;
            p_read_45_reg_3169_pp0_iter29_reg <= p_read_45_reg_3169_pp0_iter28_reg;
            p_read_45_reg_3169_pp0_iter2_reg <= p_read_45_reg_3169_pp0_iter1_reg;
            p_read_45_reg_3169_pp0_iter30_reg <= p_read_45_reg_3169_pp0_iter29_reg;
            p_read_45_reg_3169_pp0_iter31_reg <= p_read_45_reg_3169_pp0_iter30_reg;
            p_read_45_reg_3169_pp0_iter32_reg <= p_read_45_reg_3169_pp0_iter31_reg;
            p_read_45_reg_3169_pp0_iter33_reg <= p_read_45_reg_3169_pp0_iter32_reg;
            p_read_45_reg_3169_pp0_iter34_reg <= p_read_45_reg_3169_pp0_iter33_reg;
            p_read_45_reg_3169_pp0_iter35_reg <= p_read_45_reg_3169_pp0_iter34_reg;
            p_read_45_reg_3169_pp0_iter36_reg <= p_read_45_reg_3169_pp0_iter35_reg;
            p_read_45_reg_3169_pp0_iter37_reg <= p_read_45_reg_3169_pp0_iter36_reg;
            p_read_45_reg_3169_pp0_iter38_reg <= p_read_45_reg_3169_pp0_iter37_reg;
            p_read_45_reg_3169_pp0_iter39_reg <= p_read_45_reg_3169_pp0_iter38_reg;
            p_read_45_reg_3169_pp0_iter3_reg <= p_read_45_reg_3169_pp0_iter2_reg;
            p_read_45_reg_3169_pp0_iter40_reg <= p_read_45_reg_3169_pp0_iter39_reg;
            p_read_45_reg_3169_pp0_iter41_reg <= p_read_45_reg_3169_pp0_iter40_reg;
            p_read_45_reg_3169_pp0_iter42_reg <= p_read_45_reg_3169_pp0_iter41_reg;
            p_read_45_reg_3169_pp0_iter43_reg <= p_read_45_reg_3169_pp0_iter42_reg;
            p_read_45_reg_3169_pp0_iter44_reg <= p_read_45_reg_3169_pp0_iter43_reg;
            p_read_45_reg_3169_pp0_iter45_reg <= p_read_45_reg_3169_pp0_iter44_reg;
            p_read_45_reg_3169_pp0_iter46_reg <= p_read_45_reg_3169_pp0_iter45_reg;
            p_read_45_reg_3169_pp0_iter47_reg <= p_read_45_reg_3169_pp0_iter46_reg;
            p_read_45_reg_3169_pp0_iter48_reg <= p_read_45_reg_3169_pp0_iter47_reg;
            p_read_45_reg_3169_pp0_iter49_reg <= p_read_45_reg_3169_pp0_iter48_reg;
            p_read_45_reg_3169_pp0_iter4_reg <= p_read_45_reg_3169_pp0_iter3_reg;
            p_read_45_reg_3169_pp0_iter50_reg <= p_read_45_reg_3169_pp0_iter49_reg;
            p_read_45_reg_3169_pp0_iter51_reg <= p_read_45_reg_3169_pp0_iter50_reg;
            p_read_45_reg_3169_pp0_iter52_reg <= p_read_45_reg_3169_pp0_iter51_reg;
            p_read_45_reg_3169_pp0_iter53_reg <= p_read_45_reg_3169_pp0_iter52_reg;
            p_read_45_reg_3169_pp0_iter54_reg <= p_read_45_reg_3169_pp0_iter53_reg;
            p_read_45_reg_3169_pp0_iter55_reg <= p_read_45_reg_3169_pp0_iter54_reg;
            p_read_45_reg_3169_pp0_iter56_reg <= p_read_45_reg_3169_pp0_iter55_reg;
            p_read_45_reg_3169_pp0_iter57_reg <= p_read_45_reg_3169_pp0_iter56_reg;
            p_read_45_reg_3169_pp0_iter58_reg <= p_read_45_reg_3169_pp0_iter57_reg;
            p_read_45_reg_3169_pp0_iter59_reg <= p_read_45_reg_3169_pp0_iter58_reg;
            p_read_45_reg_3169_pp0_iter5_reg <= p_read_45_reg_3169_pp0_iter4_reg;
            p_read_45_reg_3169_pp0_iter60_reg <= p_read_45_reg_3169_pp0_iter59_reg;
            p_read_45_reg_3169_pp0_iter61_reg <= p_read_45_reg_3169_pp0_iter60_reg;
            p_read_45_reg_3169_pp0_iter62_reg <= p_read_45_reg_3169_pp0_iter61_reg;
            p_read_45_reg_3169_pp0_iter63_reg <= p_read_45_reg_3169_pp0_iter62_reg;
            p_read_45_reg_3169_pp0_iter64_reg <= p_read_45_reg_3169_pp0_iter63_reg;
            p_read_45_reg_3169_pp0_iter65_reg <= p_read_45_reg_3169_pp0_iter64_reg;
            p_read_45_reg_3169_pp0_iter66_reg <= p_read_45_reg_3169_pp0_iter65_reg;
            p_read_45_reg_3169_pp0_iter67_reg <= p_read_45_reg_3169_pp0_iter66_reg;
            p_read_45_reg_3169_pp0_iter68_reg <= p_read_45_reg_3169_pp0_iter67_reg;
            p_read_45_reg_3169_pp0_iter69_reg <= p_read_45_reg_3169_pp0_iter68_reg;
            p_read_45_reg_3169_pp0_iter6_reg <= p_read_45_reg_3169_pp0_iter5_reg;
            p_read_45_reg_3169_pp0_iter70_reg <= p_read_45_reg_3169_pp0_iter69_reg;
            p_read_45_reg_3169_pp0_iter71_reg <= p_read_45_reg_3169_pp0_iter70_reg;
            p_read_45_reg_3169_pp0_iter72_reg <= p_read_45_reg_3169_pp0_iter71_reg;
            p_read_45_reg_3169_pp0_iter73_reg <= p_read_45_reg_3169_pp0_iter72_reg;
            p_read_45_reg_3169_pp0_iter74_reg <= p_read_45_reg_3169_pp0_iter73_reg;
            p_read_45_reg_3169_pp0_iter75_reg <= p_read_45_reg_3169_pp0_iter74_reg;
            p_read_45_reg_3169_pp0_iter76_reg <= p_read_45_reg_3169_pp0_iter75_reg;
            p_read_45_reg_3169_pp0_iter7_reg <= p_read_45_reg_3169_pp0_iter6_reg;
            p_read_45_reg_3169_pp0_iter8_reg <= p_read_45_reg_3169_pp0_iter7_reg;
            p_read_45_reg_3169_pp0_iter9_reg <= p_read_45_reg_3169_pp0_iter8_reg;
            p_read_46_reg_3174 <= p_read18_int_reg;
            p_read_46_reg_3174_pp0_iter10_reg <= p_read_46_reg_3174_pp0_iter9_reg;
            p_read_46_reg_3174_pp0_iter11_reg <= p_read_46_reg_3174_pp0_iter10_reg;
            p_read_46_reg_3174_pp0_iter12_reg <= p_read_46_reg_3174_pp0_iter11_reg;
            p_read_46_reg_3174_pp0_iter13_reg <= p_read_46_reg_3174_pp0_iter12_reg;
            p_read_46_reg_3174_pp0_iter14_reg <= p_read_46_reg_3174_pp0_iter13_reg;
            p_read_46_reg_3174_pp0_iter15_reg <= p_read_46_reg_3174_pp0_iter14_reg;
            p_read_46_reg_3174_pp0_iter16_reg <= p_read_46_reg_3174_pp0_iter15_reg;
            p_read_46_reg_3174_pp0_iter17_reg <= p_read_46_reg_3174_pp0_iter16_reg;
            p_read_46_reg_3174_pp0_iter18_reg <= p_read_46_reg_3174_pp0_iter17_reg;
            p_read_46_reg_3174_pp0_iter19_reg <= p_read_46_reg_3174_pp0_iter18_reg;
            p_read_46_reg_3174_pp0_iter1_reg <= p_read_46_reg_3174;
            p_read_46_reg_3174_pp0_iter20_reg <= p_read_46_reg_3174_pp0_iter19_reg;
            p_read_46_reg_3174_pp0_iter21_reg <= p_read_46_reg_3174_pp0_iter20_reg;
            p_read_46_reg_3174_pp0_iter22_reg <= p_read_46_reg_3174_pp0_iter21_reg;
            p_read_46_reg_3174_pp0_iter23_reg <= p_read_46_reg_3174_pp0_iter22_reg;
            p_read_46_reg_3174_pp0_iter24_reg <= p_read_46_reg_3174_pp0_iter23_reg;
            p_read_46_reg_3174_pp0_iter25_reg <= p_read_46_reg_3174_pp0_iter24_reg;
            p_read_46_reg_3174_pp0_iter26_reg <= p_read_46_reg_3174_pp0_iter25_reg;
            p_read_46_reg_3174_pp0_iter27_reg <= p_read_46_reg_3174_pp0_iter26_reg;
            p_read_46_reg_3174_pp0_iter28_reg <= p_read_46_reg_3174_pp0_iter27_reg;
            p_read_46_reg_3174_pp0_iter29_reg <= p_read_46_reg_3174_pp0_iter28_reg;
            p_read_46_reg_3174_pp0_iter2_reg <= p_read_46_reg_3174_pp0_iter1_reg;
            p_read_46_reg_3174_pp0_iter30_reg <= p_read_46_reg_3174_pp0_iter29_reg;
            p_read_46_reg_3174_pp0_iter31_reg <= p_read_46_reg_3174_pp0_iter30_reg;
            p_read_46_reg_3174_pp0_iter32_reg <= p_read_46_reg_3174_pp0_iter31_reg;
            p_read_46_reg_3174_pp0_iter33_reg <= p_read_46_reg_3174_pp0_iter32_reg;
            p_read_46_reg_3174_pp0_iter34_reg <= p_read_46_reg_3174_pp0_iter33_reg;
            p_read_46_reg_3174_pp0_iter35_reg <= p_read_46_reg_3174_pp0_iter34_reg;
            p_read_46_reg_3174_pp0_iter36_reg <= p_read_46_reg_3174_pp0_iter35_reg;
            p_read_46_reg_3174_pp0_iter37_reg <= p_read_46_reg_3174_pp0_iter36_reg;
            p_read_46_reg_3174_pp0_iter38_reg <= p_read_46_reg_3174_pp0_iter37_reg;
            p_read_46_reg_3174_pp0_iter39_reg <= p_read_46_reg_3174_pp0_iter38_reg;
            p_read_46_reg_3174_pp0_iter3_reg <= p_read_46_reg_3174_pp0_iter2_reg;
            p_read_46_reg_3174_pp0_iter40_reg <= p_read_46_reg_3174_pp0_iter39_reg;
            p_read_46_reg_3174_pp0_iter41_reg <= p_read_46_reg_3174_pp0_iter40_reg;
            p_read_46_reg_3174_pp0_iter42_reg <= p_read_46_reg_3174_pp0_iter41_reg;
            p_read_46_reg_3174_pp0_iter43_reg <= p_read_46_reg_3174_pp0_iter42_reg;
            p_read_46_reg_3174_pp0_iter44_reg <= p_read_46_reg_3174_pp0_iter43_reg;
            p_read_46_reg_3174_pp0_iter45_reg <= p_read_46_reg_3174_pp0_iter44_reg;
            p_read_46_reg_3174_pp0_iter46_reg <= p_read_46_reg_3174_pp0_iter45_reg;
            p_read_46_reg_3174_pp0_iter47_reg <= p_read_46_reg_3174_pp0_iter46_reg;
            p_read_46_reg_3174_pp0_iter48_reg <= p_read_46_reg_3174_pp0_iter47_reg;
            p_read_46_reg_3174_pp0_iter49_reg <= p_read_46_reg_3174_pp0_iter48_reg;
            p_read_46_reg_3174_pp0_iter4_reg <= p_read_46_reg_3174_pp0_iter3_reg;
            p_read_46_reg_3174_pp0_iter50_reg <= p_read_46_reg_3174_pp0_iter49_reg;
            p_read_46_reg_3174_pp0_iter51_reg <= p_read_46_reg_3174_pp0_iter50_reg;
            p_read_46_reg_3174_pp0_iter52_reg <= p_read_46_reg_3174_pp0_iter51_reg;
            p_read_46_reg_3174_pp0_iter53_reg <= p_read_46_reg_3174_pp0_iter52_reg;
            p_read_46_reg_3174_pp0_iter54_reg <= p_read_46_reg_3174_pp0_iter53_reg;
            p_read_46_reg_3174_pp0_iter55_reg <= p_read_46_reg_3174_pp0_iter54_reg;
            p_read_46_reg_3174_pp0_iter56_reg <= p_read_46_reg_3174_pp0_iter55_reg;
            p_read_46_reg_3174_pp0_iter57_reg <= p_read_46_reg_3174_pp0_iter56_reg;
            p_read_46_reg_3174_pp0_iter58_reg <= p_read_46_reg_3174_pp0_iter57_reg;
            p_read_46_reg_3174_pp0_iter59_reg <= p_read_46_reg_3174_pp0_iter58_reg;
            p_read_46_reg_3174_pp0_iter5_reg <= p_read_46_reg_3174_pp0_iter4_reg;
            p_read_46_reg_3174_pp0_iter60_reg <= p_read_46_reg_3174_pp0_iter59_reg;
            p_read_46_reg_3174_pp0_iter61_reg <= p_read_46_reg_3174_pp0_iter60_reg;
            p_read_46_reg_3174_pp0_iter62_reg <= p_read_46_reg_3174_pp0_iter61_reg;
            p_read_46_reg_3174_pp0_iter63_reg <= p_read_46_reg_3174_pp0_iter62_reg;
            p_read_46_reg_3174_pp0_iter64_reg <= p_read_46_reg_3174_pp0_iter63_reg;
            p_read_46_reg_3174_pp0_iter65_reg <= p_read_46_reg_3174_pp0_iter64_reg;
            p_read_46_reg_3174_pp0_iter66_reg <= p_read_46_reg_3174_pp0_iter65_reg;
            p_read_46_reg_3174_pp0_iter67_reg <= p_read_46_reg_3174_pp0_iter66_reg;
            p_read_46_reg_3174_pp0_iter68_reg <= p_read_46_reg_3174_pp0_iter67_reg;
            p_read_46_reg_3174_pp0_iter69_reg <= p_read_46_reg_3174_pp0_iter68_reg;
            p_read_46_reg_3174_pp0_iter6_reg <= p_read_46_reg_3174_pp0_iter5_reg;
            p_read_46_reg_3174_pp0_iter70_reg <= p_read_46_reg_3174_pp0_iter69_reg;
            p_read_46_reg_3174_pp0_iter71_reg <= p_read_46_reg_3174_pp0_iter70_reg;
            p_read_46_reg_3174_pp0_iter72_reg <= p_read_46_reg_3174_pp0_iter71_reg;
            p_read_46_reg_3174_pp0_iter73_reg <= p_read_46_reg_3174_pp0_iter72_reg;
            p_read_46_reg_3174_pp0_iter74_reg <= p_read_46_reg_3174_pp0_iter73_reg;
            p_read_46_reg_3174_pp0_iter75_reg <= p_read_46_reg_3174_pp0_iter74_reg;
            p_read_46_reg_3174_pp0_iter76_reg <= p_read_46_reg_3174_pp0_iter75_reg;
            p_read_46_reg_3174_pp0_iter7_reg <= p_read_46_reg_3174_pp0_iter6_reg;
            p_read_46_reg_3174_pp0_iter8_reg <= p_read_46_reg_3174_pp0_iter7_reg;
            p_read_46_reg_3174_pp0_iter9_reg <= p_read_46_reg_3174_pp0_iter8_reg;
            p_read_47_reg_3179 <= p_read17_int_reg;
            p_read_47_reg_3179_pp0_iter10_reg <= p_read_47_reg_3179_pp0_iter9_reg;
            p_read_47_reg_3179_pp0_iter11_reg <= p_read_47_reg_3179_pp0_iter10_reg;
            p_read_47_reg_3179_pp0_iter12_reg <= p_read_47_reg_3179_pp0_iter11_reg;
            p_read_47_reg_3179_pp0_iter13_reg <= p_read_47_reg_3179_pp0_iter12_reg;
            p_read_47_reg_3179_pp0_iter14_reg <= p_read_47_reg_3179_pp0_iter13_reg;
            p_read_47_reg_3179_pp0_iter15_reg <= p_read_47_reg_3179_pp0_iter14_reg;
            p_read_47_reg_3179_pp0_iter16_reg <= p_read_47_reg_3179_pp0_iter15_reg;
            p_read_47_reg_3179_pp0_iter17_reg <= p_read_47_reg_3179_pp0_iter16_reg;
            p_read_47_reg_3179_pp0_iter18_reg <= p_read_47_reg_3179_pp0_iter17_reg;
            p_read_47_reg_3179_pp0_iter19_reg <= p_read_47_reg_3179_pp0_iter18_reg;
            p_read_47_reg_3179_pp0_iter1_reg <= p_read_47_reg_3179;
            p_read_47_reg_3179_pp0_iter20_reg <= p_read_47_reg_3179_pp0_iter19_reg;
            p_read_47_reg_3179_pp0_iter21_reg <= p_read_47_reg_3179_pp0_iter20_reg;
            p_read_47_reg_3179_pp0_iter22_reg <= p_read_47_reg_3179_pp0_iter21_reg;
            p_read_47_reg_3179_pp0_iter23_reg <= p_read_47_reg_3179_pp0_iter22_reg;
            p_read_47_reg_3179_pp0_iter24_reg <= p_read_47_reg_3179_pp0_iter23_reg;
            p_read_47_reg_3179_pp0_iter25_reg <= p_read_47_reg_3179_pp0_iter24_reg;
            p_read_47_reg_3179_pp0_iter26_reg <= p_read_47_reg_3179_pp0_iter25_reg;
            p_read_47_reg_3179_pp0_iter27_reg <= p_read_47_reg_3179_pp0_iter26_reg;
            p_read_47_reg_3179_pp0_iter28_reg <= p_read_47_reg_3179_pp0_iter27_reg;
            p_read_47_reg_3179_pp0_iter29_reg <= p_read_47_reg_3179_pp0_iter28_reg;
            p_read_47_reg_3179_pp0_iter2_reg <= p_read_47_reg_3179_pp0_iter1_reg;
            p_read_47_reg_3179_pp0_iter30_reg <= p_read_47_reg_3179_pp0_iter29_reg;
            p_read_47_reg_3179_pp0_iter31_reg <= p_read_47_reg_3179_pp0_iter30_reg;
            p_read_47_reg_3179_pp0_iter32_reg <= p_read_47_reg_3179_pp0_iter31_reg;
            p_read_47_reg_3179_pp0_iter33_reg <= p_read_47_reg_3179_pp0_iter32_reg;
            p_read_47_reg_3179_pp0_iter34_reg <= p_read_47_reg_3179_pp0_iter33_reg;
            p_read_47_reg_3179_pp0_iter35_reg <= p_read_47_reg_3179_pp0_iter34_reg;
            p_read_47_reg_3179_pp0_iter36_reg <= p_read_47_reg_3179_pp0_iter35_reg;
            p_read_47_reg_3179_pp0_iter37_reg <= p_read_47_reg_3179_pp0_iter36_reg;
            p_read_47_reg_3179_pp0_iter38_reg <= p_read_47_reg_3179_pp0_iter37_reg;
            p_read_47_reg_3179_pp0_iter39_reg <= p_read_47_reg_3179_pp0_iter38_reg;
            p_read_47_reg_3179_pp0_iter3_reg <= p_read_47_reg_3179_pp0_iter2_reg;
            p_read_47_reg_3179_pp0_iter40_reg <= p_read_47_reg_3179_pp0_iter39_reg;
            p_read_47_reg_3179_pp0_iter41_reg <= p_read_47_reg_3179_pp0_iter40_reg;
            p_read_47_reg_3179_pp0_iter42_reg <= p_read_47_reg_3179_pp0_iter41_reg;
            p_read_47_reg_3179_pp0_iter43_reg <= p_read_47_reg_3179_pp0_iter42_reg;
            p_read_47_reg_3179_pp0_iter44_reg <= p_read_47_reg_3179_pp0_iter43_reg;
            p_read_47_reg_3179_pp0_iter45_reg <= p_read_47_reg_3179_pp0_iter44_reg;
            p_read_47_reg_3179_pp0_iter46_reg <= p_read_47_reg_3179_pp0_iter45_reg;
            p_read_47_reg_3179_pp0_iter47_reg <= p_read_47_reg_3179_pp0_iter46_reg;
            p_read_47_reg_3179_pp0_iter48_reg <= p_read_47_reg_3179_pp0_iter47_reg;
            p_read_47_reg_3179_pp0_iter49_reg <= p_read_47_reg_3179_pp0_iter48_reg;
            p_read_47_reg_3179_pp0_iter4_reg <= p_read_47_reg_3179_pp0_iter3_reg;
            p_read_47_reg_3179_pp0_iter50_reg <= p_read_47_reg_3179_pp0_iter49_reg;
            p_read_47_reg_3179_pp0_iter51_reg <= p_read_47_reg_3179_pp0_iter50_reg;
            p_read_47_reg_3179_pp0_iter52_reg <= p_read_47_reg_3179_pp0_iter51_reg;
            p_read_47_reg_3179_pp0_iter53_reg <= p_read_47_reg_3179_pp0_iter52_reg;
            p_read_47_reg_3179_pp0_iter54_reg <= p_read_47_reg_3179_pp0_iter53_reg;
            p_read_47_reg_3179_pp0_iter55_reg <= p_read_47_reg_3179_pp0_iter54_reg;
            p_read_47_reg_3179_pp0_iter56_reg <= p_read_47_reg_3179_pp0_iter55_reg;
            p_read_47_reg_3179_pp0_iter57_reg <= p_read_47_reg_3179_pp0_iter56_reg;
            p_read_47_reg_3179_pp0_iter58_reg <= p_read_47_reg_3179_pp0_iter57_reg;
            p_read_47_reg_3179_pp0_iter59_reg <= p_read_47_reg_3179_pp0_iter58_reg;
            p_read_47_reg_3179_pp0_iter5_reg <= p_read_47_reg_3179_pp0_iter4_reg;
            p_read_47_reg_3179_pp0_iter60_reg <= p_read_47_reg_3179_pp0_iter59_reg;
            p_read_47_reg_3179_pp0_iter61_reg <= p_read_47_reg_3179_pp0_iter60_reg;
            p_read_47_reg_3179_pp0_iter62_reg <= p_read_47_reg_3179_pp0_iter61_reg;
            p_read_47_reg_3179_pp0_iter63_reg <= p_read_47_reg_3179_pp0_iter62_reg;
            p_read_47_reg_3179_pp0_iter64_reg <= p_read_47_reg_3179_pp0_iter63_reg;
            p_read_47_reg_3179_pp0_iter65_reg <= p_read_47_reg_3179_pp0_iter64_reg;
            p_read_47_reg_3179_pp0_iter66_reg <= p_read_47_reg_3179_pp0_iter65_reg;
            p_read_47_reg_3179_pp0_iter67_reg <= p_read_47_reg_3179_pp0_iter66_reg;
            p_read_47_reg_3179_pp0_iter68_reg <= p_read_47_reg_3179_pp0_iter67_reg;
            p_read_47_reg_3179_pp0_iter69_reg <= p_read_47_reg_3179_pp0_iter68_reg;
            p_read_47_reg_3179_pp0_iter6_reg <= p_read_47_reg_3179_pp0_iter5_reg;
            p_read_47_reg_3179_pp0_iter70_reg <= p_read_47_reg_3179_pp0_iter69_reg;
            p_read_47_reg_3179_pp0_iter71_reg <= p_read_47_reg_3179_pp0_iter70_reg;
            p_read_47_reg_3179_pp0_iter72_reg <= p_read_47_reg_3179_pp0_iter71_reg;
            p_read_47_reg_3179_pp0_iter73_reg <= p_read_47_reg_3179_pp0_iter72_reg;
            p_read_47_reg_3179_pp0_iter74_reg <= p_read_47_reg_3179_pp0_iter73_reg;
            p_read_47_reg_3179_pp0_iter75_reg <= p_read_47_reg_3179_pp0_iter74_reg;
            p_read_47_reg_3179_pp0_iter76_reg <= p_read_47_reg_3179_pp0_iter75_reg;
            p_read_47_reg_3179_pp0_iter7_reg <= p_read_47_reg_3179_pp0_iter6_reg;
            p_read_47_reg_3179_pp0_iter8_reg <= p_read_47_reg_3179_pp0_iter7_reg;
            p_read_47_reg_3179_pp0_iter9_reg <= p_read_47_reg_3179_pp0_iter8_reg;
            p_read_48_reg_3184 <= p_read16_int_reg;
            p_read_48_reg_3184_pp0_iter10_reg <= p_read_48_reg_3184_pp0_iter9_reg;
            p_read_48_reg_3184_pp0_iter11_reg <= p_read_48_reg_3184_pp0_iter10_reg;
            p_read_48_reg_3184_pp0_iter12_reg <= p_read_48_reg_3184_pp0_iter11_reg;
            p_read_48_reg_3184_pp0_iter13_reg <= p_read_48_reg_3184_pp0_iter12_reg;
            p_read_48_reg_3184_pp0_iter14_reg <= p_read_48_reg_3184_pp0_iter13_reg;
            p_read_48_reg_3184_pp0_iter15_reg <= p_read_48_reg_3184_pp0_iter14_reg;
            p_read_48_reg_3184_pp0_iter16_reg <= p_read_48_reg_3184_pp0_iter15_reg;
            p_read_48_reg_3184_pp0_iter17_reg <= p_read_48_reg_3184_pp0_iter16_reg;
            p_read_48_reg_3184_pp0_iter18_reg <= p_read_48_reg_3184_pp0_iter17_reg;
            p_read_48_reg_3184_pp0_iter19_reg <= p_read_48_reg_3184_pp0_iter18_reg;
            p_read_48_reg_3184_pp0_iter1_reg <= p_read_48_reg_3184;
            p_read_48_reg_3184_pp0_iter20_reg <= p_read_48_reg_3184_pp0_iter19_reg;
            p_read_48_reg_3184_pp0_iter21_reg <= p_read_48_reg_3184_pp0_iter20_reg;
            p_read_48_reg_3184_pp0_iter22_reg <= p_read_48_reg_3184_pp0_iter21_reg;
            p_read_48_reg_3184_pp0_iter23_reg <= p_read_48_reg_3184_pp0_iter22_reg;
            p_read_48_reg_3184_pp0_iter24_reg <= p_read_48_reg_3184_pp0_iter23_reg;
            p_read_48_reg_3184_pp0_iter25_reg <= p_read_48_reg_3184_pp0_iter24_reg;
            p_read_48_reg_3184_pp0_iter26_reg <= p_read_48_reg_3184_pp0_iter25_reg;
            p_read_48_reg_3184_pp0_iter27_reg <= p_read_48_reg_3184_pp0_iter26_reg;
            p_read_48_reg_3184_pp0_iter28_reg <= p_read_48_reg_3184_pp0_iter27_reg;
            p_read_48_reg_3184_pp0_iter29_reg <= p_read_48_reg_3184_pp0_iter28_reg;
            p_read_48_reg_3184_pp0_iter2_reg <= p_read_48_reg_3184_pp0_iter1_reg;
            p_read_48_reg_3184_pp0_iter30_reg <= p_read_48_reg_3184_pp0_iter29_reg;
            p_read_48_reg_3184_pp0_iter31_reg <= p_read_48_reg_3184_pp0_iter30_reg;
            p_read_48_reg_3184_pp0_iter32_reg <= p_read_48_reg_3184_pp0_iter31_reg;
            p_read_48_reg_3184_pp0_iter33_reg <= p_read_48_reg_3184_pp0_iter32_reg;
            p_read_48_reg_3184_pp0_iter34_reg <= p_read_48_reg_3184_pp0_iter33_reg;
            p_read_48_reg_3184_pp0_iter35_reg <= p_read_48_reg_3184_pp0_iter34_reg;
            p_read_48_reg_3184_pp0_iter36_reg <= p_read_48_reg_3184_pp0_iter35_reg;
            p_read_48_reg_3184_pp0_iter37_reg <= p_read_48_reg_3184_pp0_iter36_reg;
            p_read_48_reg_3184_pp0_iter38_reg <= p_read_48_reg_3184_pp0_iter37_reg;
            p_read_48_reg_3184_pp0_iter39_reg <= p_read_48_reg_3184_pp0_iter38_reg;
            p_read_48_reg_3184_pp0_iter3_reg <= p_read_48_reg_3184_pp0_iter2_reg;
            p_read_48_reg_3184_pp0_iter40_reg <= p_read_48_reg_3184_pp0_iter39_reg;
            p_read_48_reg_3184_pp0_iter41_reg <= p_read_48_reg_3184_pp0_iter40_reg;
            p_read_48_reg_3184_pp0_iter42_reg <= p_read_48_reg_3184_pp0_iter41_reg;
            p_read_48_reg_3184_pp0_iter43_reg <= p_read_48_reg_3184_pp0_iter42_reg;
            p_read_48_reg_3184_pp0_iter44_reg <= p_read_48_reg_3184_pp0_iter43_reg;
            p_read_48_reg_3184_pp0_iter45_reg <= p_read_48_reg_3184_pp0_iter44_reg;
            p_read_48_reg_3184_pp0_iter46_reg <= p_read_48_reg_3184_pp0_iter45_reg;
            p_read_48_reg_3184_pp0_iter47_reg <= p_read_48_reg_3184_pp0_iter46_reg;
            p_read_48_reg_3184_pp0_iter48_reg <= p_read_48_reg_3184_pp0_iter47_reg;
            p_read_48_reg_3184_pp0_iter49_reg <= p_read_48_reg_3184_pp0_iter48_reg;
            p_read_48_reg_3184_pp0_iter4_reg <= p_read_48_reg_3184_pp0_iter3_reg;
            p_read_48_reg_3184_pp0_iter50_reg <= p_read_48_reg_3184_pp0_iter49_reg;
            p_read_48_reg_3184_pp0_iter51_reg <= p_read_48_reg_3184_pp0_iter50_reg;
            p_read_48_reg_3184_pp0_iter52_reg <= p_read_48_reg_3184_pp0_iter51_reg;
            p_read_48_reg_3184_pp0_iter53_reg <= p_read_48_reg_3184_pp0_iter52_reg;
            p_read_48_reg_3184_pp0_iter54_reg <= p_read_48_reg_3184_pp0_iter53_reg;
            p_read_48_reg_3184_pp0_iter55_reg <= p_read_48_reg_3184_pp0_iter54_reg;
            p_read_48_reg_3184_pp0_iter56_reg <= p_read_48_reg_3184_pp0_iter55_reg;
            p_read_48_reg_3184_pp0_iter57_reg <= p_read_48_reg_3184_pp0_iter56_reg;
            p_read_48_reg_3184_pp0_iter58_reg <= p_read_48_reg_3184_pp0_iter57_reg;
            p_read_48_reg_3184_pp0_iter59_reg <= p_read_48_reg_3184_pp0_iter58_reg;
            p_read_48_reg_3184_pp0_iter5_reg <= p_read_48_reg_3184_pp0_iter4_reg;
            p_read_48_reg_3184_pp0_iter60_reg <= p_read_48_reg_3184_pp0_iter59_reg;
            p_read_48_reg_3184_pp0_iter61_reg <= p_read_48_reg_3184_pp0_iter60_reg;
            p_read_48_reg_3184_pp0_iter62_reg <= p_read_48_reg_3184_pp0_iter61_reg;
            p_read_48_reg_3184_pp0_iter63_reg <= p_read_48_reg_3184_pp0_iter62_reg;
            p_read_48_reg_3184_pp0_iter64_reg <= p_read_48_reg_3184_pp0_iter63_reg;
            p_read_48_reg_3184_pp0_iter65_reg <= p_read_48_reg_3184_pp0_iter64_reg;
            p_read_48_reg_3184_pp0_iter66_reg <= p_read_48_reg_3184_pp0_iter65_reg;
            p_read_48_reg_3184_pp0_iter67_reg <= p_read_48_reg_3184_pp0_iter66_reg;
            p_read_48_reg_3184_pp0_iter68_reg <= p_read_48_reg_3184_pp0_iter67_reg;
            p_read_48_reg_3184_pp0_iter69_reg <= p_read_48_reg_3184_pp0_iter68_reg;
            p_read_48_reg_3184_pp0_iter6_reg <= p_read_48_reg_3184_pp0_iter5_reg;
            p_read_48_reg_3184_pp0_iter70_reg <= p_read_48_reg_3184_pp0_iter69_reg;
            p_read_48_reg_3184_pp0_iter71_reg <= p_read_48_reg_3184_pp0_iter70_reg;
            p_read_48_reg_3184_pp0_iter72_reg <= p_read_48_reg_3184_pp0_iter71_reg;
            p_read_48_reg_3184_pp0_iter73_reg <= p_read_48_reg_3184_pp0_iter72_reg;
            p_read_48_reg_3184_pp0_iter74_reg <= p_read_48_reg_3184_pp0_iter73_reg;
            p_read_48_reg_3184_pp0_iter75_reg <= p_read_48_reg_3184_pp0_iter74_reg;
            p_read_48_reg_3184_pp0_iter76_reg <= p_read_48_reg_3184_pp0_iter75_reg;
            p_read_48_reg_3184_pp0_iter7_reg <= p_read_48_reg_3184_pp0_iter6_reg;
            p_read_48_reg_3184_pp0_iter8_reg <= p_read_48_reg_3184_pp0_iter7_reg;
            p_read_48_reg_3184_pp0_iter9_reg <= p_read_48_reg_3184_pp0_iter8_reg;
            p_read_49_reg_3189 <= p_read15_int_reg;
            p_read_49_reg_3189_pp0_iter10_reg <= p_read_49_reg_3189_pp0_iter9_reg;
            p_read_49_reg_3189_pp0_iter11_reg <= p_read_49_reg_3189_pp0_iter10_reg;
            p_read_49_reg_3189_pp0_iter12_reg <= p_read_49_reg_3189_pp0_iter11_reg;
            p_read_49_reg_3189_pp0_iter13_reg <= p_read_49_reg_3189_pp0_iter12_reg;
            p_read_49_reg_3189_pp0_iter14_reg <= p_read_49_reg_3189_pp0_iter13_reg;
            p_read_49_reg_3189_pp0_iter15_reg <= p_read_49_reg_3189_pp0_iter14_reg;
            p_read_49_reg_3189_pp0_iter16_reg <= p_read_49_reg_3189_pp0_iter15_reg;
            p_read_49_reg_3189_pp0_iter17_reg <= p_read_49_reg_3189_pp0_iter16_reg;
            p_read_49_reg_3189_pp0_iter18_reg <= p_read_49_reg_3189_pp0_iter17_reg;
            p_read_49_reg_3189_pp0_iter19_reg <= p_read_49_reg_3189_pp0_iter18_reg;
            p_read_49_reg_3189_pp0_iter1_reg <= p_read_49_reg_3189;
            p_read_49_reg_3189_pp0_iter20_reg <= p_read_49_reg_3189_pp0_iter19_reg;
            p_read_49_reg_3189_pp0_iter21_reg <= p_read_49_reg_3189_pp0_iter20_reg;
            p_read_49_reg_3189_pp0_iter22_reg <= p_read_49_reg_3189_pp0_iter21_reg;
            p_read_49_reg_3189_pp0_iter23_reg <= p_read_49_reg_3189_pp0_iter22_reg;
            p_read_49_reg_3189_pp0_iter24_reg <= p_read_49_reg_3189_pp0_iter23_reg;
            p_read_49_reg_3189_pp0_iter25_reg <= p_read_49_reg_3189_pp0_iter24_reg;
            p_read_49_reg_3189_pp0_iter26_reg <= p_read_49_reg_3189_pp0_iter25_reg;
            p_read_49_reg_3189_pp0_iter27_reg <= p_read_49_reg_3189_pp0_iter26_reg;
            p_read_49_reg_3189_pp0_iter28_reg <= p_read_49_reg_3189_pp0_iter27_reg;
            p_read_49_reg_3189_pp0_iter29_reg <= p_read_49_reg_3189_pp0_iter28_reg;
            p_read_49_reg_3189_pp0_iter2_reg <= p_read_49_reg_3189_pp0_iter1_reg;
            p_read_49_reg_3189_pp0_iter30_reg <= p_read_49_reg_3189_pp0_iter29_reg;
            p_read_49_reg_3189_pp0_iter31_reg <= p_read_49_reg_3189_pp0_iter30_reg;
            p_read_49_reg_3189_pp0_iter32_reg <= p_read_49_reg_3189_pp0_iter31_reg;
            p_read_49_reg_3189_pp0_iter33_reg <= p_read_49_reg_3189_pp0_iter32_reg;
            p_read_49_reg_3189_pp0_iter34_reg <= p_read_49_reg_3189_pp0_iter33_reg;
            p_read_49_reg_3189_pp0_iter35_reg <= p_read_49_reg_3189_pp0_iter34_reg;
            p_read_49_reg_3189_pp0_iter36_reg <= p_read_49_reg_3189_pp0_iter35_reg;
            p_read_49_reg_3189_pp0_iter37_reg <= p_read_49_reg_3189_pp0_iter36_reg;
            p_read_49_reg_3189_pp0_iter38_reg <= p_read_49_reg_3189_pp0_iter37_reg;
            p_read_49_reg_3189_pp0_iter39_reg <= p_read_49_reg_3189_pp0_iter38_reg;
            p_read_49_reg_3189_pp0_iter3_reg <= p_read_49_reg_3189_pp0_iter2_reg;
            p_read_49_reg_3189_pp0_iter40_reg <= p_read_49_reg_3189_pp0_iter39_reg;
            p_read_49_reg_3189_pp0_iter41_reg <= p_read_49_reg_3189_pp0_iter40_reg;
            p_read_49_reg_3189_pp0_iter42_reg <= p_read_49_reg_3189_pp0_iter41_reg;
            p_read_49_reg_3189_pp0_iter43_reg <= p_read_49_reg_3189_pp0_iter42_reg;
            p_read_49_reg_3189_pp0_iter44_reg <= p_read_49_reg_3189_pp0_iter43_reg;
            p_read_49_reg_3189_pp0_iter45_reg <= p_read_49_reg_3189_pp0_iter44_reg;
            p_read_49_reg_3189_pp0_iter46_reg <= p_read_49_reg_3189_pp0_iter45_reg;
            p_read_49_reg_3189_pp0_iter47_reg <= p_read_49_reg_3189_pp0_iter46_reg;
            p_read_49_reg_3189_pp0_iter48_reg <= p_read_49_reg_3189_pp0_iter47_reg;
            p_read_49_reg_3189_pp0_iter49_reg <= p_read_49_reg_3189_pp0_iter48_reg;
            p_read_49_reg_3189_pp0_iter4_reg <= p_read_49_reg_3189_pp0_iter3_reg;
            p_read_49_reg_3189_pp0_iter50_reg <= p_read_49_reg_3189_pp0_iter49_reg;
            p_read_49_reg_3189_pp0_iter51_reg <= p_read_49_reg_3189_pp0_iter50_reg;
            p_read_49_reg_3189_pp0_iter52_reg <= p_read_49_reg_3189_pp0_iter51_reg;
            p_read_49_reg_3189_pp0_iter53_reg <= p_read_49_reg_3189_pp0_iter52_reg;
            p_read_49_reg_3189_pp0_iter54_reg <= p_read_49_reg_3189_pp0_iter53_reg;
            p_read_49_reg_3189_pp0_iter55_reg <= p_read_49_reg_3189_pp0_iter54_reg;
            p_read_49_reg_3189_pp0_iter56_reg <= p_read_49_reg_3189_pp0_iter55_reg;
            p_read_49_reg_3189_pp0_iter57_reg <= p_read_49_reg_3189_pp0_iter56_reg;
            p_read_49_reg_3189_pp0_iter58_reg <= p_read_49_reg_3189_pp0_iter57_reg;
            p_read_49_reg_3189_pp0_iter59_reg <= p_read_49_reg_3189_pp0_iter58_reg;
            p_read_49_reg_3189_pp0_iter5_reg <= p_read_49_reg_3189_pp0_iter4_reg;
            p_read_49_reg_3189_pp0_iter60_reg <= p_read_49_reg_3189_pp0_iter59_reg;
            p_read_49_reg_3189_pp0_iter61_reg <= p_read_49_reg_3189_pp0_iter60_reg;
            p_read_49_reg_3189_pp0_iter62_reg <= p_read_49_reg_3189_pp0_iter61_reg;
            p_read_49_reg_3189_pp0_iter63_reg <= p_read_49_reg_3189_pp0_iter62_reg;
            p_read_49_reg_3189_pp0_iter64_reg <= p_read_49_reg_3189_pp0_iter63_reg;
            p_read_49_reg_3189_pp0_iter65_reg <= p_read_49_reg_3189_pp0_iter64_reg;
            p_read_49_reg_3189_pp0_iter66_reg <= p_read_49_reg_3189_pp0_iter65_reg;
            p_read_49_reg_3189_pp0_iter67_reg <= p_read_49_reg_3189_pp0_iter66_reg;
            p_read_49_reg_3189_pp0_iter68_reg <= p_read_49_reg_3189_pp0_iter67_reg;
            p_read_49_reg_3189_pp0_iter69_reg <= p_read_49_reg_3189_pp0_iter68_reg;
            p_read_49_reg_3189_pp0_iter6_reg <= p_read_49_reg_3189_pp0_iter5_reg;
            p_read_49_reg_3189_pp0_iter70_reg <= p_read_49_reg_3189_pp0_iter69_reg;
            p_read_49_reg_3189_pp0_iter71_reg <= p_read_49_reg_3189_pp0_iter70_reg;
            p_read_49_reg_3189_pp0_iter72_reg <= p_read_49_reg_3189_pp0_iter71_reg;
            p_read_49_reg_3189_pp0_iter73_reg <= p_read_49_reg_3189_pp0_iter72_reg;
            p_read_49_reg_3189_pp0_iter74_reg <= p_read_49_reg_3189_pp0_iter73_reg;
            p_read_49_reg_3189_pp0_iter75_reg <= p_read_49_reg_3189_pp0_iter74_reg;
            p_read_49_reg_3189_pp0_iter76_reg <= p_read_49_reg_3189_pp0_iter75_reg;
            p_read_49_reg_3189_pp0_iter7_reg <= p_read_49_reg_3189_pp0_iter6_reg;
            p_read_49_reg_3189_pp0_iter8_reg <= p_read_49_reg_3189_pp0_iter7_reg;
            p_read_49_reg_3189_pp0_iter9_reg <= p_read_49_reg_3189_pp0_iter8_reg;
            p_read_50_reg_3194 <= p_read14_int_reg;
            p_read_50_reg_3194_pp0_iter10_reg <= p_read_50_reg_3194_pp0_iter9_reg;
            p_read_50_reg_3194_pp0_iter11_reg <= p_read_50_reg_3194_pp0_iter10_reg;
            p_read_50_reg_3194_pp0_iter12_reg <= p_read_50_reg_3194_pp0_iter11_reg;
            p_read_50_reg_3194_pp0_iter13_reg <= p_read_50_reg_3194_pp0_iter12_reg;
            p_read_50_reg_3194_pp0_iter14_reg <= p_read_50_reg_3194_pp0_iter13_reg;
            p_read_50_reg_3194_pp0_iter15_reg <= p_read_50_reg_3194_pp0_iter14_reg;
            p_read_50_reg_3194_pp0_iter16_reg <= p_read_50_reg_3194_pp0_iter15_reg;
            p_read_50_reg_3194_pp0_iter17_reg <= p_read_50_reg_3194_pp0_iter16_reg;
            p_read_50_reg_3194_pp0_iter18_reg <= p_read_50_reg_3194_pp0_iter17_reg;
            p_read_50_reg_3194_pp0_iter19_reg <= p_read_50_reg_3194_pp0_iter18_reg;
            p_read_50_reg_3194_pp0_iter1_reg <= p_read_50_reg_3194;
            p_read_50_reg_3194_pp0_iter20_reg <= p_read_50_reg_3194_pp0_iter19_reg;
            p_read_50_reg_3194_pp0_iter21_reg <= p_read_50_reg_3194_pp0_iter20_reg;
            p_read_50_reg_3194_pp0_iter22_reg <= p_read_50_reg_3194_pp0_iter21_reg;
            p_read_50_reg_3194_pp0_iter23_reg <= p_read_50_reg_3194_pp0_iter22_reg;
            p_read_50_reg_3194_pp0_iter24_reg <= p_read_50_reg_3194_pp0_iter23_reg;
            p_read_50_reg_3194_pp0_iter25_reg <= p_read_50_reg_3194_pp0_iter24_reg;
            p_read_50_reg_3194_pp0_iter26_reg <= p_read_50_reg_3194_pp0_iter25_reg;
            p_read_50_reg_3194_pp0_iter27_reg <= p_read_50_reg_3194_pp0_iter26_reg;
            p_read_50_reg_3194_pp0_iter28_reg <= p_read_50_reg_3194_pp0_iter27_reg;
            p_read_50_reg_3194_pp0_iter29_reg <= p_read_50_reg_3194_pp0_iter28_reg;
            p_read_50_reg_3194_pp0_iter2_reg <= p_read_50_reg_3194_pp0_iter1_reg;
            p_read_50_reg_3194_pp0_iter30_reg <= p_read_50_reg_3194_pp0_iter29_reg;
            p_read_50_reg_3194_pp0_iter31_reg <= p_read_50_reg_3194_pp0_iter30_reg;
            p_read_50_reg_3194_pp0_iter32_reg <= p_read_50_reg_3194_pp0_iter31_reg;
            p_read_50_reg_3194_pp0_iter33_reg <= p_read_50_reg_3194_pp0_iter32_reg;
            p_read_50_reg_3194_pp0_iter34_reg <= p_read_50_reg_3194_pp0_iter33_reg;
            p_read_50_reg_3194_pp0_iter35_reg <= p_read_50_reg_3194_pp0_iter34_reg;
            p_read_50_reg_3194_pp0_iter36_reg <= p_read_50_reg_3194_pp0_iter35_reg;
            p_read_50_reg_3194_pp0_iter37_reg <= p_read_50_reg_3194_pp0_iter36_reg;
            p_read_50_reg_3194_pp0_iter38_reg <= p_read_50_reg_3194_pp0_iter37_reg;
            p_read_50_reg_3194_pp0_iter39_reg <= p_read_50_reg_3194_pp0_iter38_reg;
            p_read_50_reg_3194_pp0_iter3_reg <= p_read_50_reg_3194_pp0_iter2_reg;
            p_read_50_reg_3194_pp0_iter40_reg <= p_read_50_reg_3194_pp0_iter39_reg;
            p_read_50_reg_3194_pp0_iter41_reg <= p_read_50_reg_3194_pp0_iter40_reg;
            p_read_50_reg_3194_pp0_iter42_reg <= p_read_50_reg_3194_pp0_iter41_reg;
            p_read_50_reg_3194_pp0_iter43_reg <= p_read_50_reg_3194_pp0_iter42_reg;
            p_read_50_reg_3194_pp0_iter44_reg <= p_read_50_reg_3194_pp0_iter43_reg;
            p_read_50_reg_3194_pp0_iter45_reg <= p_read_50_reg_3194_pp0_iter44_reg;
            p_read_50_reg_3194_pp0_iter46_reg <= p_read_50_reg_3194_pp0_iter45_reg;
            p_read_50_reg_3194_pp0_iter47_reg <= p_read_50_reg_3194_pp0_iter46_reg;
            p_read_50_reg_3194_pp0_iter48_reg <= p_read_50_reg_3194_pp0_iter47_reg;
            p_read_50_reg_3194_pp0_iter49_reg <= p_read_50_reg_3194_pp0_iter48_reg;
            p_read_50_reg_3194_pp0_iter4_reg <= p_read_50_reg_3194_pp0_iter3_reg;
            p_read_50_reg_3194_pp0_iter50_reg <= p_read_50_reg_3194_pp0_iter49_reg;
            p_read_50_reg_3194_pp0_iter51_reg <= p_read_50_reg_3194_pp0_iter50_reg;
            p_read_50_reg_3194_pp0_iter52_reg <= p_read_50_reg_3194_pp0_iter51_reg;
            p_read_50_reg_3194_pp0_iter53_reg <= p_read_50_reg_3194_pp0_iter52_reg;
            p_read_50_reg_3194_pp0_iter54_reg <= p_read_50_reg_3194_pp0_iter53_reg;
            p_read_50_reg_3194_pp0_iter55_reg <= p_read_50_reg_3194_pp0_iter54_reg;
            p_read_50_reg_3194_pp0_iter56_reg <= p_read_50_reg_3194_pp0_iter55_reg;
            p_read_50_reg_3194_pp0_iter57_reg <= p_read_50_reg_3194_pp0_iter56_reg;
            p_read_50_reg_3194_pp0_iter58_reg <= p_read_50_reg_3194_pp0_iter57_reg;
            p_read_50_reg_3194_pp0_iter59_reg <= p_read_50_reg_3194_pp0_iter58_reg;
            p_read_50_reg_3194_pp0_iter5_reg <= p_read_50_reg_3194_pp0_iter4_reg;
            p_read_50_reg_3194_pp0_iter60_reg <= p_read_50_reg_3194_pp0_iter59_reg;
            p_read_50_reg_3194_pp0_iter61_reg <= p_read_50_reg_3194_pp0_iter60_reg;
            p_read_50_reg_3194_pp0_iter62_reg <= p_read_50_reg_3194_pp0_iter61_reg;
            p_read_50_reg_3194_pp0_iter63_reg <= p_read_50_reg_3194_pp0_iter62_reg;
            p_read_50_reg_3194_pp0_iter64_reg <= p_read_50_reg_3194_pp0_iter63_reg;
            p_read_50_reg_3194_pp0_iter65_reg <= p_read_50_reg_3194_pp0_iter64_reg;
            p_read_50_reg_3194_pp0_iter66_reg <= p_read_50_reg_3194_pp0_iter65_reg;
            p_read_50_reg_3194_pp0_iter67_reg <= p_read_50_reg_3194_pp0_iter66_reg;
            p_read_50_reg_3194_pp0_iter68_reg <= p_read_50_reg_3194_pp0_iter67_reg;
            p_read_50_reg_3194_pp0_iter69_reg <= p_read_50_reg_3194_pp0_iter68_reg;
            p_read_50_reg_3194_pp0_iter6_reg <= p_read_50_reg_3194_pp0_iter5_reg;
            p_read_50_reg_3194_pp0_iter70_reg <= p_read_50_reg_3194_pp0_iter69_reg;
            p_read_50_reg_3194_pp0_iter71_reg <= p_read_50_reg_3194_pp0_iter70_reg;
            p_read_50_reg_3194_pp0_iter72_reg <= p_read_50_reg_3194_pp0_iter71_reg;
            p_read_50_reg_3194_pp0_iter73_reg <= p_read_50_reg_3194_pp0_iter72_reg;
            p_read_50_reg_3194_pp0_iter74_reg <= p_read_50_reg_3194_pp0_iter73_reg;
            p_read_50_reg_3194_pp0_iter75_reg <= p_read_50_reg_3194_pp0_iter74_reg;
            p_read_50_reg_3194_pp0_iter76_reg <= p_read_50_reg_3194_pp0_iter75_reg;
            p_read_50_reg_3194_pp0_iter7_reg <= p_read_50_reg_3194_pp0_iter6_reg;
            p_read_50_reg_3194_pp0_iter8_reg <= p_read_50_reg_3194_pp0_iter7_reg;
            p_read_50_reg_3194_pp0_iter9_reg <= p_read_50_reg_3194_pp0_iter8_reg;
            p_read_51_reg_3199 <= p_read13_int_reg;
            p_read_51_reg_3199_pp0_iter10_reg <= p_read_51_reg_3199_pp0_iter9_reg;
            p_read_51_reg_3199_pp0_iter11_reg <= p_read_51_reg_3199_pp0_iter10_reg;
            p_read_51_reg_3199_pp0_iter12_reg <= p_read_51_reg_3199_pp0_iter11_reg;
            p_read_51_reg_3199_pp0_iter13_reg <= p_read_51_reg_3199_pp0_iter12_reg;
            p_read_51_reg_3199_pp0_iter14_reg <= p_read_51_reg_3199_pp0_iter13_reg;
            p_read_51_reg_3199_pp0_iter15_reg <= p_read_51_reg_3199_pp0_iter14_reg;
            p_read_51_reg_3199_pp0_iter16_reg <= p_read_51_reg_3199_pp0_iter15_reg;
            p_read_51_reg_3199_pp0_iter17_reg <= p_read_51_reg_3199_pp0_iter16_reg;
            p_read_51_reg_3199_pp0_iter18_reg <= p_read_51_reg_3199_pp0_iter17_reg;
            p_read_51_reg_3199_pp0_iter19_reg <= p_read_51_reg_3199_pp0_iter18_reg;
            p_read_51_reg_3199_pp0_iter1_reg <= p_read_51_reg_3199;
            p_read_51_reg_3199_pp0_iter20_reg <= p_read_51_reg_3199_pp0_iter19_reg;
            p_read_51_reg_3199_pp0_iter21_reg <= p_read_51_reg_3199_pp0_iter20_reg;
            p_read_51_reg_3199_pp0_iter22_reg <= p_read_51_reg_3199_pp0_iter21_reg;
            p_read_51_reg_3199_pp0_iter23_reg <= p_read_51_reg_3199_pp0_iter22_reg;
            p_read_51_reg_3199_pp0_iter24_reg <= p_read_51_reg_3199_pp0_iter23_reg;
            p_read_51_reg_3199_pp0_iter25_reg <= p_read_51_reg_3199_pp0_iter24_reg;
            p_read_51_reg_3199_pp0_iter26_reg <= p_read_51_reg_3199_pp0_iter25_reg;
            p_read_51_reg_3199_pp0_iter27_reg <= p_read_51_reg_3199_pp0_iter26_reg;
            p_read_51_reg_3199_pp0_iter28_reg <= p_read_51_reg_3199_pp0_iter27_reg;
            p_read_51_reg_3199_pp0_iter29_reg <= p_read_51_reg_3199_pp0_iter28_reg;
            p_read_51_reg_3199_pp0_iter2_reg <= p_read_51_reg_3199_pp0_iter1_reg;
            p_read_51_reg_3199_pp0_iter30_reg <= p_read_51_reg_3199_pp0_iter29_reg;
            p_read_51_reg_3199_pp0_iter31_reg <= p_read_51_reg_3199_pp0_iter30_reg;
            p_read_51_reg_3199_pp0_iter32_reg <= p_read_51_reg_3199_pp0_iter31_reg;
            p_read_51_reg_3199_pp0_iter33_reg <= p_read_51_reg_3199_pp0_iter32_reg;
            p_read_51_reg_3199_pp0_iter34_reg <= p_read_51_reg_3199_pp0_iter33_reg;
            p_read_51_reg_3199_pp0_iter35_reg <= p_read_51_reg_3199_pp0_iter34_reg;
            p_read_51_reg_3199_pp0_iter36_reg <= p_read_51_reg_3199_pp0_iter35_reg;
            p_read_51_reg_3199_pp0_iter37_reg <= p_read_51_reg_3199_pp0_iter36_reg;
            p_read_51_reg_3199_pp0_iter38_reg <= p_read_51_reg_3199_pp0_iter37_reg;
            p_read_51_reg_3199_pp0_iter39_reg <= p_read_51_reg_3199_pp0_iter38_reg;
            p_read_51_reg_3199_pp0_iter3_reg <= p_read_51_reg_3199_pp0_iter2_reg;
            p_read_51_reg_3199_pp0_iter40_reg <= p_read_51_reg_3199_pp0_iter39_reg;
            p_read_51_reg_3199_pp0_iter41_reg <= p_read_51_reg_3199_pp0_iter40_reg;
            p_read_51_reg_3199_pp0_iter42_reg <= p_read_51_reg_3199_pp0_iter41_reg;
            p_read_51_reg_3199_pp0_iter43_reg <= p_read_51_reg_3199_pp0_iter42_reg;
            p_read_51_reg_3199_pp0_iter44_reg <= p_read_51_reg_3199_pp0_iter43_reg;
            p_read_51_reg_3199_pp0_iter45_reg <= p_read_51_reg_3199_pp0_iter44_reg;
            p_read_51_reg_3199_pp0_iter46_reg <= p_read_51_reg_3199_pp0_iter45_reg;
            p_read_51_reg_3199_pp0_iter47_reg <= p_read_51_reg_3199_pp0_iter46_reg;
            p_read_51_reg_3199_pp0_iter48_reg <= p_read_51_reg_3199_pp0_iter47_reg;
            p_read_51_reg_3199_pp0_iter49_reg <= p_read_51_reg_3199_pp0_iter48_reg;
            p_read_51_reg_3199_pp0_iter4_reg <= p_read_51_reg_3199_pp0_iter3_reg;
            p_read_51_reg_3199_pp0_iter50_reg <= p_read_51_reg_3199_pp0_iter49_reg;
            p_read_51_reg_3199_pp0_iter51_reg <= p_read_51_reg_3199_pp0_iter50_reg;
            p_read_51_reg_3199_pp0_iter52_reg <= p_read_51_reg_3199_pp0_iter51_reg;
            p_read_51_reg_3199_pp0_iter53_reg <= p_read_51_reg_3199_pp0_iter52_reg;
            p_read_51_reg_3199_pp0_iter54_reg <= p_read_51_reg_3199_pp0_iter53_reg;
            p_read_51_reg_3199_pp0_iter55_reg <= p_read_51_reg_3199_pp0_iter54_reg;
            p_read_51_reg_3199_pp0_iter56_reg <= p_read_51_reg_3199_pp0_iter55_reg;
            p_read_51_reg_3199_pp0_iter57_reg <= p_read_51_reg_3199_pp0_iter56_reg;
            p_read_51_reg_3199_pp0_iter58_reg <= p_read_51_reg_3199_pp0_iter57_reg;
            p_read_51_reg_3199_pp0_iter59_reg <= p_read_51_reg_3199_pp0_iter58_reg;
            p_read_51_reg_3199_pp0_iter5_reg <= p_read_51_reg_3199_pp0_iter4_reg;
            p_read_51_reg_3199_pp0_iter60_reg <= p_read_51_reg_3199_pp0_iter59_reg;
            p_read_51_reg_3199_pp0_iter61_reg <= p_read_51_reg_3199_pp0_iter60_reg;
            p_read_51_reg_3199_pp0_iter62_reg <= p_read_51_reg_3199_pp0_iter61_reg;
            p_read_51_reg_3199_pp0_iter63_reg <= p_read_51_reg_3199_pp0_iter62_reg;
            p_read_51_reg_3199_pp0_iter64_reg <= p_read_51_reg_3199_pp0_iter63_reg;
            p_read_51_reg_3199_pp0_iter65_reg <= p_read_51_reg_3199_pp0_iter64_reg;
            p_read_51_reg_3199_pp0_iter66_reg <= p_read_51_reg_3199_pp0_iter65_reg;
            p_read_51_reg_3199_pp0_iter67_reg <= p_read_51_reg_3199_pp0_iter66_reg;
            p_read_51_reg_3199_pp0_iter68_reg <= p_read_51_reg_3199_pp0_iter67_reg;
            p_read_51_reg_3199_pp0_iter69_reg <= p_read_51_reg_3199_pp0_iter68_reg;
            p_read_51_reg_3199_pp0_iter6_reg <= p_read_51_reg_3199_pp0_iter5_reg;
            p_read_51_reg_3199_pp0_iter70_reg <= p_read_51_reg_3199_pp0_iter69_reg;
            p_read_51_reg_3199_pp0_iter71_reg <= p_read_51_reg_3199_pp0_iter70_reg;
            p_read_51_reg_3199_pp0_iter72_reg <= p_read_51_reg_3199_pp0_iter71_reg;
            p_read_51_reg_3199_pp0_iter73_reg <= p_read_51_reg_3199_pp0_iter72_reg;
            p_read_51_reg_3199_pp0_iter74_reg <= p_read_51_reg_3199_pp0_iter73_reg;
            p_read_51_reg_3199_pp0_iter75_reg <= p_read_51_reg_3199_pp0_iter74_reg;
            p_read_51_reg_3199_pp0_iter76_reg <= p_read_51_reg_3199_pp0_iter75_reg;
            p_read_51_reg_3199_pp0_iter7_reg <= p_read_51_reg_3199_pp0_iter6_reg;
            p_read_51_reg_3199_pp0_iter8_reg <= p_read_51_reg_3199_pp0_iter7_reg;
            p_read_51_reg_3199_pp0_iter9_reg <= p_read_51_reg_3199_pp0_iter8_reg;
            p_read_52_reg_3204 <= p_read12_int_reg;
            p_read_52_reg_3204_pp0_iter10_reg <= p_read_52_reg_3204_pp0_iter9_reg;
            p_read_52_reg_3204_pp0_iter11_reg <= p_read_52_reg_3204_pp0_iter10_reg;
            p_read_52_reg_3204_pp0_iter12_reg <= p_read_52_reg_3204_pp0_iter11_reg;
            p_read_52_reg_3204_pp0_iter13_reg <= p_read_52_reg_3204_pp0_iter12_reg;
            p_read_52_reg_3204_pp0_iter14_reg <= p_read_52_reg_3204_pp0_iter13_reg;
            p_read_52_reg_3204_pp0_iter15_reg <= p_read_52_reg_3204_pp0_iter14_reg;
            p_read_52_reg_3204_pp0_iter16_reg <= p_read_52_reg_3204_pp0_iter15_reg;
            p_read_52_reg_3204_pp0_iter17_reg <= p_read_52_reg_3204_pp0_iter16_reg;
            p_read_52_reg_3204_pp0_iter18_reg <= p_read_52_reg_3204_pp0_iter17_reg;
            p_read_52_reg_3204_pp0_iter19_reg <= p_read_52_reg_3204_pp0_iter18_reg;
            p_read_52_reg_3204_pp0_iter1_reg <= p_read_52_reg_3204;
            p_read_52_reg_3204_pp0_iter20_reg <= p_read_52_reg_3204_pp0_iter19_reg;
            p_read_52_reg_3204_pp0_iter21_reg <= p_read_52_reg_3204_pp0_iter20_reg;
            p_read_52_reg_3204_pp0_iter22_reg <= p_read_52_reg_3204_pp0_iter21_reg;
            p_read_52_reg_3204_pp0_iter23_reg <= p_read_52_reg_3204_pp0_iter22_reg;
            p_read_52_reg_3204_pp0_iter24_reg <= p_read_52_reg_3204_pp0_iter23_reg;
            p_read_52_reg_3204_pp0_iter25_reg <= p_read_52_reg_3204_pp0_iter24_reg;
            p_read_52_reg_3204_pp0_iter26_reg <= p_read_52_reg_3204_pp0_iter25_reg;
            p_read_52_reg_3204_pp0_iter27_reg <= p_read_52_reg_3204_pp0_iter26_reg;
            p_read_52_reg_3204_pp0_iter28_reg <= p_read_52_reg_3204_pp0_iter27_reg;
            p_read_52_reg_3204_pp0_iter29_reg <= p_read_52_reg_3204_pp0_iter28_reg;
            p_read_52_reg_3204_pp0_iter2_reg <= p_read_52_reg_3204_pp0_iter1_reg;
            p_read_52_reg_3204_pp0_iter30_reg <= p_read_52_reg_3204_pp0_iter29_reg;
            p_read_52_reg_3204_pp0_iter31_reg <= p_read_52_reg_3204_pp0_iter30_reg;
            p_read_52_reg_3204_pp0_iter32_reg <= p_read_52_reg_3204_pp0_iter31_reg;
            p_read_52_reg_3204_pp0_iter33_reg <= p_read_52_reg_3204_pp0_iter32_reg;
            p_read_52_reg_3204_pp0_iter34_reg <= p_read_52_reg_3204_pp0_iter33_reg;
            p_read_52_reg_3204_pp0_iter35_reg <= p_read_52_reg_3204_pp0_iter34_reg;
            p_read_52_reg_3204_pp0_iter36_reg <= p_read_52_reg_3204_pp0_iter35_reg;
            p_read_52_reg_3204_pp0_iter37_reg <= p_read_52_reg_3204_pp0_iter36_reg;
            p_read_52_reg_3204_pp0_iter38_reg <= p_read_52_reg_3204_pp0_iter37_reg;
            p_read_52_reg_3204_pp0_iter39_reg <= p_read_52_reg_3204_pp0_iter38_reg;
            p_read_52_reg_3204_pp0_iter3_reg <= p_read_52_reg_3204_pp0_iter2_reg;
            p_read_52_reg_3204_pp0_iter40_reg <= p_read_52_reg_3204_pp0_iter39_reg;
            p_read_52_reg_3204_pp0_iter41_reg <= p_read_52_reg_3204_pp0_iter40_reg;
            p_read_52_reg_3204_pp0_iter42_reg <= p_read_52_reg_3204_pp0_iter41_reg;
            p_read_52_reg_3204_pp0_iter43_reg <= p_read_52_reg_3204_pp0_iter42_reg;
            p_read_52_reg_3204_pp0_iter44_reg <= p_read_52_reg_3204_pp0_iter43_reg;
            p_read_52_reg_3204_pp0_iter45_reg <= p_read_52_reg_3204_pp0_iter44_reg;
            p_read_52_reg_3204_pp0_iter46_reg <= p_read_52_reg_3204_pp0_iter45_reg;
            p_read_52_reg_3204_pp0_iter47_reg <= p_read_52_reg_3204_pp0_iter46_reg;
            p_read_52_reg_3204_pp0_iter48_reg <= p_read_52_reg_3204_pp0_iter47_reg;
            p_read_52_reg_3204_pp0_iter49_reg <= p_read_52_reg_3204_pp0_iter48_reg;
            p_read_52_reg_3204_pp0_iter4_reg <= p_read_52_reg_3204_pp0_iter3_reg;
            p_read_52_reg_3204_pp0_iter50_reg <= p_read_52_reg_3204_pp0_iter49_reg;
            p_read_52_reg_3204_pp0_iter51_reg <= p_read_52_reg_3204_pp0_iter50_reg;
            p_read_52_reg_3204_pp0_iter52_reg <= p_read_52_reg_3204_pp0_iter51_reg;
            p_read_52_reg_3204_pp0_iter53_reg <= p_read_52_reg_3204_pp0_iter52_reg;
            p_read_52_reg_3204_pp0_iter54_reg <= p_read_52_reg_3204_pp0_iter53_reg;
            p_read_52_reg_3204_pp0_iter55_reg <= p_read_52_reg_3204_pp0_iter54_reg;
            p_read_52_reg_3204_pp0_iter56_reg <= p_read_52_reg_3204_pp0_iter55_reg;
            p_read_52_reg_3204_pp0_iter57_reg <= p_read_52_reg_3204_pp0_iter56_reg;
            p_read_52_reg_3204_pp0_iter58_reg <= p_read_52_reg_3204_pp0_iter57_reg;
            p_read_52_reg_3204_pp0_iter59_reg <= p_read_52_reg_3204_pp0_iter58_reg;
            p_read_52_reg_3204_pp0_iter5_reg <= p_read_52_reg_3204_pp0_iter4_reg;
            p_read_52_reg_3204_pp0_iter60_reg <= p_read_52_reg_3204_pp0_iter59_reg;
            p_read_52_reg_3204_pp0_iter61_reg <= p_read_52_reg_3204_pp0_iter60_reg;
            p_read_52_reg_3204_pp0_iter62_reg <= p_read_52_reg_3204_pp0_iter61_reg;
            p_read_52_reg_3204_pp0_iter63_reg <= p_read_52_reg_3204_pp0_iter62_reg;
            p_read_52_reg_3204_pp0_iter64_reg <= p_read_52_reg_3204_pp0_iter63_reg;
            p_read_52_reg_3204_pp0_iter65_reg <= p_read_52_reg_3204_pp0_iter64_reg;
            p_read_52_reg_3204_pp0_iter66_reg <= p_read_52_reg_3204_pp0_iter65_reg;
            p_read_52_reg_3204_pp0_iter67_reg <= p_read_52_reg_3204_pp0_iter66_reg;
            p_read_52_reg_3204_pp0_iter68_reg <= p_read_52_reg_3204_pp0_iter67_reg;
            p_read_52_reg_3204_pp0_iter69_reg <= p_read_52_reg_3204_pp0_iter68_reg;
            p_read_52_reg_3204_pp0_iter6_reg <= p_read_52_reg_3204_pp0_iter5_reg;
            p_read_52_reg_3204_pp0_iter70_reg <= p_read_52_reg_3204_pp0_iter69_reg;
            p_read_52_reg_3204_pp0_iter71_reg <= p_read_52_reg_3204_pp0_iter70_reg;
            p_read_52_reg_3204_pp0_iter72_reg <= p_read_52_reg_3204_pp0_iter71_reg;
            p_read_52_reg_3204_pp0_iter73_reg <= p_read_52_reg_3204_pp0_iter72_reg;
            p_read_52_reg_3204_pp0_iter74_reg <= p_read_52_reg_3204_pp0_iter73_reg;
            p_read_52_reg_3204_pp0_iter75_reg <= p_read_52_reg_3204_pp0_iter74_reg;
            p_read_52_reg_3204_pp0_iter76_reg <= p_read_52_reg_3204_pp0_iter75_reg;
            p_read_52_reg_3204_pp0_iter7_reg <= p_read_52_reg_3204_pp0_iter6_reg;
            p_read_52_reg_3204_pp0_iter8_reg <= p_read_52_reg_3204_pp0_iter7_reg;
            p_read_52_reg_3204_pp0_iter9_reg <= p_read_52_reg_3204_pp0_iter8_reg;
            p_read_53_reg_3209 <= p_read11_int_reg;
            p_read_53_reg_3209_pp0_iter10_reg <= p_read_53_reg_3209_pp0_iter9_reg;
            p_read_53_reg_3209_pp0_iter11_reg <= p_read_53_reg_3209_pp0_iter10_reg;
            p_read_53_reg_3209_pp0_iter12_reg <= p_read_53_reg_3209_pp0_iter11_reg;
            p_read_53_reg_3209_pp0_iter13_reg <= p_read_53_reg_3209_pp0_iter12_reg;
            p_read_53_reg_3209_pp0_iter14_reg <= p_read_53_reg_3209_pp0_iter13_reg;
            p_read_53_reg_3209_pp0_iter15_reg <= p_read_53_reg_3209_pp0_iter14_reg;
            p_read_53_reg_3209_pp0_iter16_reg <= p_read_53_reg_3209_pp0_iter15_reg;
            p_read_53_reg_3209_pp0_iter17_reg <= p_read_53_reg_3209_pp0_iter16_reg;
            p_read_53_reg_3209_pp0_iter18_reg <= p_read_53_reg_3209_pp0_iter17_reg;
            p_read_53_reg_3209_pp0_iter19_reg <= p_read_53_reg_3209_pp0_iter18_reg;
            p_read_53_reg_3209_pp0_iter1_reg <= p_read_53_reg_3209;
            p_read_53_reg_3209_pp0_iter20_reg <= p_read_53_reg_3209_pp0_iter19_reg;
            p_read_53_reg_3209_pp0_iter21_reg <= p_read_53_reg_3209_pp0_iter20_reg;
            p_read_53_reg_3209_pp0_iter22_reg <= p_read_53_reg_3209_pp0_iter21_reg;
            p_read_53_reg_3209_pp0_iter23_reg <= p_read_53_reg_3209_pp0_iter22_reg;
            p_read_53_reg_3209_pp0_iter24_reg <= p_read_53_reg_3209_pp0_iter23_reg;
            p_read_53_reg_3209_pp0_iter25_reg <= p_read_53_reg_3209_pp0_iter24_reg;
            p_read_53_reg_3209_pp0_iter26_reg <= p_read_53_reg_3209_pp0_iter25_reg;
            p_read_53_reg_3209_pp0_iter27_reg <= p_read_53_reg_3209_pp0_iter26_reg;
            p_read_53_reg_3209_pp0_iter28_reg <= p_read_53_reg_3209_pp0_iter27_reg;
            p_read_53_reg_3209_pp0_iter29_reg <= p_read_53_reg_3209_pp0_iter28_reg;
            p_read_53_reg_3209_pp0_iter2_reg <= p_read_53_reg_3209_pp0_iter1_reg;
            p_read_53_reg_3209_pp0_iter30_reg <= p_read_53_reg_3209_pp0_iter29_reg;
            p_read_53_reg_3209_pp0_iter31_reg <= p_read_53_reg_3209_pp0_iter30_reg;
            p_read_53_reg_3209_pp0_iter32_reg <= p_read_53_reg_3209_pp0_iter31_reg;
            p_read_53_reg_3209_pp0_iter33_reg <= p_read_53_reg_3209_pp0_iter32_reg;
            p_read_53_reg_3209_pp0_iter34_reg <= p_read_53_reg_3209_pp0_iter33_reg;
            p_read_53_reg_3209_pp0_iter35_reg <= p_read_53_reg_3209_pp0_iter34_reg;
            p_read_53_reg_3209_pp0_iter36_reg <= p_read_53_reg_3209_pp0_iter35_reg;
            p_read_53_reg_3209_pp0_iter37_reg <= p_read_53_reg_3209_pp0_iter36_reg;
            p_read_53_reg_3209_pp0_iter38_reg <= p_read_53_reg_3209_pp0_iter37_reg;
            p_read_53_reg_3209_pp0_iter39_reg <= p_read_53_reg_3209_pp0_iter38_reg;
            p_read_53_reg_3209_pp0_iter3_reg <= p_read_53_reg_3209_pp0_iter2_reg;
            p_read_53_reg_3209_pp0_iter40_reg <= p_read_53_reg_3209_pp0_iter39_reg;
            p_read_53_reg_3209_pp0_iter41_reg <= p_read_53_reg_3209_pp0_iter40_reg;
            p_read_53_reg_3209_pp0_iter42_reg <= p_read_53_reg_3209_pp0_iter41_reg;
            p_read_53_reg_3209_pp0_iter43_reg <= p_read_53_reg_3209_pp0_iter42_reg;
            p_read_53_reg_3209_pp0_iter44_reg <= p_read_53_reg_3209_pp0_iter43_reg;
            p_read_53_reg_3209_pp0_iter45_reg <= p_read_53_reg_3209_pp0_iter44_reg;
            p_read_53_reg_3209_pp0_iter46_reg <= p_read_53_reg_3209_pp0_iter45_reg;
            p_read_53_reg_3209_pp0_iter47_reg <= p_read_53_reg_3209_pp0_iter46_reg;
            p_read_53_reg_3209_pp0_iter48_reg <= p_read_53_reg_3209_pp0_iter47_reg;
            p_read_53_reg_3209_pp0_iter49_reg <= p_read_53_reg_3209_pp0_iter48_reg;
            p_read_53_reg_3209_pp0_iter4_reg <= p_read_53_reg_3209_pp0_iter3_reg;
            p_read_53_reg_3209_pp0_iter50_reg <= p_read_53_reg_3209_pp0_iter49_reg;
            p_read_53_reg_3209_pp0_iter51_reg <= p_read_53_reg_3209_pp0_iter50_reg;
            p_read_53_reg_3209_pp0_iter52_reg <= p_read_53_reg_3209_pp0_iter51_reg;
            p_read_53_reg_3209_pp0_iter53_reg <= p_read_53_reg_3209_pp0_iter52_reg;
            p_read_53_reg_3209_pp0_iter54_reg <= p_read_53_reg_3209_pp0_iter53_reg;
            p_read_53_reg_3209_pp0_iter55_reg <= p_read_53_reg_3209_pp0_iter54_reg;
            p_read_53_reg_3209_pp0_iter56_reg <= p_read_53_reg_3209_pp0_iter55_reg;
            p_read_53_reg_3209_pp0_iter57_reg <= p_read_53_reg_3209_pp0_iter56_reg;
            p_read_53_reg_3209_pp0_iter58_reg <= p_read_53_reg_3209_pp0_iter57_reg;
            p_read_53_reg_3209_pp0_iter59_reg <= p_read_53_reg_3209_pp0_iter58_reg;
            p_read_53_reg_3209_pp0_iter5_reg <= p_read_53_reg_3209_pp0_iter4_reg;
            p_read_53_reg_3209_pp0_iter60_reg <= p_read_53_reg_3209_pp0_iter59_reg;
            p_read_53_reg_3209_pp0_iter61_reg <= p_read_53_reg_3209_pp0_iter60_reg;
            p_read_53_reg_3209_pp0_iter62_reg <= p_read_53_reg_3209_pp0_iter61_reg;
            p_read_53_reg_3209_pp0_iter63_reg <= p_read_53_reg_3209_pp0_iter62_reg;
            p_read_53_reg_3209_pp0_iter64_reg <= p_read_53_reg_3209_pp0_iter63_reg;
            p_read_53_reg_3209_pp0_iter65_reg <= p_read_53_reg_3209_pp0_iter64_reg;
            p_read_53_reg_3209_pp0_iter66_reg <= p_read_53_reg_3209_pp0_iter65_reg;
            p_read_53_reg_3209_pp0_iter67_reg <= p_read_53_reg_3209_pp0_iter66_reg;
            p_read_53_reg_3209_pp0_iter68_reg <= p_read_53_reg_3209_pp0_iter67_reg;
            p_read_53_reg_3209_pp0_iter69_reg <= p_read_53_reg_3209_pp0_iter68_reg;
            p_read_53_reg_3209_pp0_iter6_reg <= p_read_53_reg_3209_pp0_iter5_reg;
            p_read_53_reg_3209_pp0_iter70_reg <= p_read_53_reg_3209_pp0_iter69_reg;
            p_read_53_reg_3209_pp0_iter71_reg <= p_read_53_reg_3209_pp0_iter70_reg;
            p_read_53_reg_3209_pp0_iter72_reg <= p_read_53_reg_3209_pp0_iter71_reg;
            p_read_53_reg_3209_pp0_iter73_reg <= p_read_53_reg_3209_pp0_iter72_reg;
            p_read_53_reg_3209_pp0_iter74_reg <= p_read_53_reg_3209_pp0_iter73_reg;
            p_read_53_reg_3209_pp0_iter75_reg <= p_read_53_reg_3209_pp0_iter74_reg;
            p_read_53_reg_3209_pp0_iter76_reg <= p_read_53_reg_3209_pp0_iter75_reg;
            p_read_53_reg_3209_pp0_iter7_reg <= p_read_53_reg_3209_pp0_iter6_reg;
            p_read_53_reg_3209_pp0_iter8_reg <= p_read_53_reg_3209_pp0_iter7_reg;
            p_read_53_reg_3209_pp0_iter9_reg <= p_read_53_reg_3209_pp0_iter8_reg;
            p_read_54_reg_3214 <= p_read10_int_reg;
            p_read_54_reg_3214_pp0_iter10_reg <= p_read_54_reg_3214_pp0_iter9_reg;
            p_read_54_reg_3214_pp0_iter11_reg <= p_read_54_reg_3214_pp0_iter10_reg;
            p_read_54_reg_3214_pp0_iter12_reg <= p_read_54_reg_3214_pp0_iter11_reg;
            p_read_54_reg_3214_pp0_iter13_reg <= p_read_54_reg_3214_pp0_iter12_reg;
            p_read_54_reg_3214_pp0_iter14_reg <= p_read_54_reg_3214_pp0_iter13_reg;
            p_read_54_reg_3214_pp0_iter15_reg <= p_read_54_reg_3214_pp0_iter14_reg;
            p_read_54_reg_3214_pp0_iter16_reg <= p_read_54_reg_3214_pp0_iter15_reg;
            p_read_54_reg_3214_pp0_iter17_reg <= p_read_54_reg_3214_pp0_iter16_reg;
            p_read_54_reg_3214_pp0_iter18_reg <= p_read_54_reg_3214_pp0_iter17_reg;
            p_read_54_reg_3214_pp0_iter19_reg <= p_read_54_reg_3214_pp0_iter18_reg;
            p_read_54_reg_3214_pp0_iter1_reg <= p_read_54_reg_3214;
            p_read_54_reg_3214_pp0_iter20_reg <= p_read_54_reg_3214_pp0_iter19_reg;
            p_read_54_reg_3214_pp0_iter21_reg <= p_read_54_reg_3214_pp0_iter20_reg;
            p_read_54_reg_3214_pp0_iter22_reg <= p_read_54_reg_3214_pp0_iter21_reg;
            p_read_54_reg_3214_pp0_iter23_reg <= p_read_54_reg_3214_pp0_iter22_reg;
            p_read_54_reg_3214_pp0_iter24_reg <= p_read_54_reg_3214_pp0_iter23_reg;
            p_read_54_reg_3214_pp0_iter25_reg <= p_read_54_reg_3214_pp0_iter24_reg;
            p_read_54_reg_3214_pp0_iter26_reg <= p_read_54_reg_3214_pp0_iter25_reg;
            p_read_54_reg_3214_pp0_iter27_reg <= p_read_54_reg_3214_pp0_iter26_reg;
            p_read_54_reg_3214_pp0_iter28_reg <= p_read_54_reg_3214_pp0_iter27_reg;
            p_read_54_reg_3214_pp0_iter29_reg <= p_read_54_reg_3214_pp0_iter28_reg;
            p_read_54_reg_3214_pp0_iter2_reg <= p_read_54_reg_3214_pp0_iter1_reg;
            p_read_54_reg_3214_pp0_iter30_reg <= p_read_54_reg_3214_pp0_iter29_reg;
            p_read_54_reg_3214_pp0_iter31_reg <= p_read_54_reg_3214_pp0_iter30_reg;
            p_read_54_reg_3214_pp0_iter32_reg <= p_read_54_reg_3214_pp0_iter31_reg;
            p_read_54_reg_3214_pp0_iter33_reg <= p_read_54_reg_3214_pp0_iter32_reg;
            p_read_54_reg_3214_pp0_iter34_reg <= p_read_54_reg_3214_pp0_iter33_reg;
            p_read_54_reg_3214_pp0_iter35_reg <= p_read_54_reg_3214_pp0_iter34_reg;
            p_read_54_reg_3214_pp0_iter36_reg <= p_read_54_reg_3214_pp0_iter35_reg;
            p_read_54_reg_3214_pp0_iter37_reg <= p_read_54_reg_3214_pp0_iter36_reg;
            p_read_54_reg_3214_pp0_iter38_reg <= p_read_54_reg_3214_pp0_iter37_reg;
            p_read_54_reg_3214_pp0_iter39_reg <= p_read_54_reg_3214_pp0_iter38_reg;
            p_read_54_reg_3214_pp0_iter3_reg <= p_read_54_reg_3214_pp0_iter2_reg;
            p_read_54_reg_3214_pp0_iter40_reg <= p_read_54_reg_3214_pp0_iter39_reg;
            p_read_54_reg_3214_pp0_iter41_reg <= p_read_54_reg_3214_pp0_iter40_reg;
            p_read_54_reg_3214_pp0_iter42_reg <= p_read_54_reg_3214_pp0_iter41_reg;
            p_read_54_reg_3214_pp0_iter43_reg <= p_read_54_reg_3214_pp0_iter42_reg;
            p_read_54_reg_3214_pp0_iter44_reg <= p_read_54_reg_3214_pp0_iter43_reg;
            p_read_54_reg_3214_pp0_iter45_reg <= p_read_54_reg_3214_pp0_iter44_reg;
            p_read_54_reg_3214_pp0_iter46_reg <= p_read_54_reg_3214_pp0_iter45_reg;
            p_read_54_reg_3214_pp0_iter47_reg <= p_read_54_reg_3214_pp0_iter46_reg;
            p_read_54_reg_3214_pp0_iter48_reg <= p_read_54_reg_3214_pp0_iter47_reg;
            p_read_54_reg_3214_pp0_iter49_reg <= p_read_54_reg_3214_pp0_iter48_reg;
            p_read_54_reg_3214_pp0_iter4_reg <= p_read_54_reg_3214_pp0_iter3_reg;
            p_read_54_reg_3214_pp0_iter50_reg <= p_read_54_reg_3214_pp0_iter49_reg;
            p_read_54_reg_3214_pp0_iter51_reg <= p_read_54_reg_3214_pp0_iter50_reg;
            p_read_54_reg_3214_pp0_iter52_reg <= p_read_54_reg_3214_pp0_iter51_reg;
            p_read_54_reg_3214_pp0_iter53_reg <= p_read_54_reg_3214_pp0_iter52_reg;
            p_read_54_reg_3214_pp0_iter54_reg <= p_read_54_reg_3214_pp0_iter53_reg;
            p_read_54_reg_3214_pp0_iter55_reg <= p_read_54_reg_3214_pp0_iter54_reg;
            p_read_54_reg_3214_pp0_iter56_reg <= p_read_54_reg_3214_pp0_iter55_reg;
            p_read_54_reg_3214_pp0_iter57_reg <= p_read_54_reg_3214_pp0_iter56_reg;
            p_read_54_reg_3214_pp0_iter58_reg <= p_read_54_reg_3214_pp0_iter57_reg;
            p_read_54_reg_3214_pp0_iter59_reg <= p_read_54_reg_3214_pp0_iter58_reg;
            p_read_54_reg_3214_pp0_iter5_reg <= p_read_54_reg_3214_pp0_iter4_reg;
            p_read_54_reg_3214_pp0_iter60_reg <= p_read_54_reg_3214_pp0_iter59_reg;
            p_read_54_reg_3214_pp0_iter61_reg <= p_read_54_reg_3214_pp0_iter60_reg;
            p_read_54_reg_3214_pp0_iter62_reg <= p_read_54_reg_3214_pp0_iter61_reg;
            p_read_54_reg_3214_pp0_iter63_reg <= p_read_54_reg_3214_pp0_iter62_reg;
            p_read_54_reg_3214_pp0_iter64_reg <= p_read_54_reg_3214_pp0_iter63_reg;
            p_read_54_reg_3214_pp0_iter65_reg <= p_read_54_reg_3214_pp0_iter64_reg;
            p_read_54_reg_3214_pp0_iter66_reg <= p_read_54_reg_3214_pp0_iter65_reg;
            p_read_54_reg_3214_pp0_iter67_reg <= p_read_54_reg_3214_pp0_iter66_reg;
            p_read_54_reg_3214_pp0_iter68_reg <= p_read_54_reg_3214_pp0_iter67_reg;
            p_read_54_reg_3214_pp0_iter69_reg <= p_read_54_reg_3214_pp0_iter68_reg;
            p_read_54_reg_3214_pp0_iter6_reg <= p_read_54_reg_3214_pp0_iter5_reg;
            p_read_54_reg_3214_pp0_iter70_reg <= p_read_54_reg_3214_pp0_iter69_reg;
            p_read_54_reg_3214_pp0_iter71_reg <= p_read_54_reg_3214_pp0_iter70_reg;
            p_read_54_reg_3214_pp0_iter72_reg <= p_read_54_reg_3214_pp0_iter71_reg;
            p_read_54_reg_3214_pp0_iter73_reg <= p_read_54_reg_3214_pp0_iter72_reg;
            p_read_54_reg_3214_pp0_iter74_reg <= p_read_54_reg_3214_pp0_iter73_reg;
            p_read_54_reg_3214_pp0_iter75_reg <= p_read_54_reg_3214_pp0_iter74_reg;
            p_read_54_reg_3214_pp0_iter76_reg <= p_read_54_reg_3214_pp0_iter75_reg;
            p_read_54_reg_3214_pp0_iter7_reg <= p_read_54_reg_3214_pp0_iter6_reg;
            p_read_54_reg_3214_pp0_iter8_reg <= p_read_54_reg_3214_pp0_iter7_reg;
            p_read_54_reg_3214_pp0_iter9_reg <= p_read_54_reg_3214_pp0_iter8_reg;
            p_read_55_reg_3219 <= p_read9_int_reg;
            p_read_55_reg_3219_pp0_iter10_reg <= p_read_55_reg_3219_pp0_iter9_reg;
            p_read_55_reg_3219_pp0_iter11_reg <= p_read_55_reg_3219_pp0_iter10_reg;
            p_read_55_reg_3219_pp0_iter12_reg <= p_read_55_reg_3219_pp0_iter11_reg;
            p_read_55_reg_3219_pp0_iter13_reg <= p_read_55_reg_3219_pp0_iter12_reg;
            p_read_55_reg_3219_pp0_iter14_reg <= p_read_55_reg_3219_pp0_iter13_reg;
            p_read_55_reg_3219_pp0_iter15_reg <= p_read_55_reg_3219_pp0_iter14_reg;
            p_read_55_reg_3219_pp0_iter16_reg <= p_read_55_reg_3219_pp0_iter15_reg;
            p_read_55_reg_3219_pp0_iter17_reg <= p_read_55_reg_3219_pp0_iter16_reg;
            p_read_55_reg_3219_pp0_iter18_reg <= p_read_55_reg_3219_pp0_iter17_reg;
            p_read_55_reg_3219_pp0_iter19_reg <= p_read_55_reg_3219_pp0_iter18_reg;
            p_read_55_reg_3219_pp0_iter1_reg <= p_read_55_reg_3219;
            p_read_55_reg_3219_pp0_iter20_reg <= p_read_55_reg_3219_pp0_iter19_reg;
            p_read_55_reg_3219_pp0_iter21_reg <= p_read_55_reg_3219_pp0_iter20_reg;
            p_read_55_reg_3219_pp0_iter22_reg <= p_read_55_reg_3219_pp0_iter21_reg;
            p_read_55_reg_3219_pp0_iter23_reg <= p_read_55_reg_3219_pp0_iter22_reg;
            p_read_55_reg_3219_pp0_iter24_reg <= p_read_55_reg_3219_pp0_iter23_reg;
            p_read_55_reg_3219_pp0_iter25_reg <= p_read_55_reg_3219_pp0_iter24_reg;
            p_read_55_reg_3219_pp0_iter26_reg <= p_read_55_reg_3219_pp0_iter25_reg;
            p_read_55_reg_3219_pp0_iter27_reg <= p_read_55_reg_3219_pp0_iter26_reg;
            p_read_55_reg_3219_pp0_iter28_reg <= p_read_55_reg_3219_pp0_iter27_reg;
            p_read_55_reg_3219_pp0_iter29_reg <= p_read_55_reg_3219_pp0_iter28_reg;
            p_read_55_reg_3219_pp0_iter2_reg <= p_read_55_reg_3219_pp0_iter1_reg;
            p_read_55_reg_3219_pp0_iter30_reg <= p_read_55_reg_3219_pp0_iter29_reg;
            p_read_55_reg_3219_pp0_iter31_reg <= p_read_55_reg_3219_pp0_iter30_reg;
            p_read_55_reg_3219_pp0_iter32_reg <= p_read_55_reg_3219_pp0_iter31_reg;
            p_read_55_reg_3219_pp0_iter33_reg <= p_read_55_reg_3219_pp0_iter32_reg;
            p_read_55_reg_3219_pp0_iter34_reg <= p_read_55_reg_3219_pp0_iter33_reg;
            p_read_55_reg_3219_pp0_iter35_reg <= p_read_55_reg_3219_pp0_iter34_reg;
            p_read_55_reg_3219_pp0_iter36_reg <= p_read_55_reg_3219_pp0_iter35_reg;
            p_read_55_reg_3219_pp0_iter37_reg <= p_read_55_reg_3219_pp0_iter36_reg;
            p_read_55_reg_3219_pp0_iter38_reg <= p_read_55_reg_3219_pp0_iter37_reg;
            p_read_55_reg_3219_pp0_iter39_reg <= p_read_55_reg_3219_pp0_iter38_reg;
            p_read_55_reg_3219_pp0_iter3_reg <= p_read_55_reg_3219_pp0_iter2_reg;
            p_read_55_reg_3219_pp0_iter40_reg <= p_read_55_reg_3219_pp0_iter39_reg;
            p_read_55_reg_3219_pp0_iter41_reg <= p_read_55_reg_3219_pp0_iter40_reg;
            p_read_55_reg_3219_pp0_iter42_reg <= p_read_55_reg_3219_pp0_iter41_reg;
            p_read_55_reg_3219_pp0_iter43_reg <= p_read_55_reg_3219_pp0_iter42_reg;
            p_read_55_reg_3219_pp0_iter44_reg <= p_read_55_reg_3219_pp0_iter43_reg;
            p_read_55_reg_3219_pp0_iter45_reg <= p_read_55_reg_3219_pp0_iter44_reg;
            p_read_55_reg_3219_pp0_iter46_reg <= p_read_55_reg_3219_pp0_iter45_reg;
            p_read_55_reg_3219_pp0_iter47_reg <= p_read_55_reg_3219_pp0_iter46_reg;
            p_read_55_reg_3219_pp0_iter48_reg <= p_read_55_reg_3219_pp0_iter47_reg;
            p_read_55_reg_3219_pp0_iter49_reg <= p_read_55_reg_3219_pp0_iter48_reg;
            p_read_55_reg_3219_pp0_iter4_reg <= p_read_55_reg_3219_pp0_iter3_reg;
            p_read_55_reg_3219_pp0_iter50_reg <= p_read_55_reg_3219_pp0_iter49_reg;
            p_read_55_reg_3219_pp0_iter51_reg <= p_read_55_reg_3219_pp0_iter50_reg;
            p_read_55_reg_3219_pp0_iter52_reg <= p_read_55_reg_3219_pp0_iter51_reg;
            p_read_55_reg_3219_pp0_iter53_reg <= p_read_55_reg_3219_pp0_iter52_reg;
            p_read_55_reg_3219_pp0_iter54_reg <= p_read_55_reg_3219_pp0_iter53_reg;
            p_read_55_reg_3219_pp0_iter55_reg <= p_read_55_reg_3219_pp0_iter54_reg;
            p_read_55_reg_3219_pp0_iter56_reg <= p_read_55_reg_3219_pp0_iter55_reg;
            p_read_55_reg_3219_pp0_iter57_reg <= p_read_55_reg_3219_pp0_iter56_reg;
            p_read_55_reg_3219_pp0_iter58_reg <= p_read_55_reg_3219_pp0_iter57_reg;
            p_read_55_reg_3219_pp0_iter59_reg <= p_read_55_reg_3219_pp0_iter58_reg;
            p_read_55_reg_3219_pp0_iter5_reg <= p_read_55_reg_3219_pp0_iter4_reg;
            p_read_55_reg_3219_pp0_iter60_reg <= p_read_55_reg_3219_pp0_iter59_reg;
            p_read_55_reg_3219_pp0_iter61_reg <= p_read_55_reg_3219_pp0_iter60_reg;
            p_read_55_reg_3219_pp0_iter62_reg <= p_read_55_reg_3219_pp0_iter61_reg;
            p_read_55_reg_3219_pp0_iter63_reg <= p_read_55_reg_3219_pp0_iter62_reg;
            p_read_55_reg_3219_pp0_iter64_reg <= p_read_55_reg_3219_pp0_iter63_reg;
            p_read_55_reg_3219_pp0_iter65_reg <= p_read_55_reg_3219_pp0_iter64_reg;
            p_read_55_reg_3219_pp0_iter66_reg <= p_read_55_reg_3219_pp0_iter65_reg;
            p_read_55_reg_3219_pp0_iter67_reg <= p_read_55_reg_3219_pp0_iter66_reg;
            p_read_55_reg_3219_pp0_iter68_reg <= p_read_55_reg_3219_pp0_iter67_reg;
            p_read_55_reg_3219_pp0_iter69_reg <= p_read_55_reg_3219_pp0_iter68_reg;
            p_read_55_reg_3219_pp0_iter6_reg <= p_read_55_reg_3219_pp0_iter5_reg;
            p_read_55_reg_3219_pp0_iter70_reg <= p_read_55_reg_3219_pp0_iter69_reg;
            p_read_55_reg_3219_pp0_iter71_reg <= p_read_55_reg_3219_pp0_iter70_reg;
            p_read_55_reg_3219_pp0_iter72_reg <= p_read_55_reg_3219_pp0_iter71_reg;
            p_read_55_reg_3219_pp0_iter73_reg <= p_read_55_reg_3219_pp0_iter72_reg;
            p_read_55_reg_3219_pp0_iter74_reg <= p_read_55_reg_3219_pp0_iter73_reg;
            p_read_55_reg_3219_pp0_iter75_reg <= p_read_55_reg_3219_pp0_iter74_reg;
            p_read_55_reg_3219_pp0_iter76_reg <= p_read_55_reg_3219_pp0_iter75_reg;
            p_read_55_reg_3219_pp0_iter7_reg <= p_read_55_reg_3219_pp0_iter6_reg;
            p_read_55_reg_3219_pp0_iter8_reg <= p_read_55_reg_3219_pp0_iter7_reg;
            p_read_55_reg_3219_pp0_iter9_reg <= p_read_55_reg_3219_pp0_iter8_reg;
            p_read_56_reg_3224 <= p_read8_int_reg;
            p_read_56_reg_3224_pp0_iter10_reg <= p_read_56_reg_3224_pp0_iter9_reg;
            p_read_56_reg_3224_pp0_iter11_reg <= p_read_56_reg_3224_pp0_iter10_reg;
            p_read_56_reg_3224_pp0_iter12_reg <= p_read_56_reg_3224_pp0_iter11_reg;
            p_read_56_reg_3224_pp0_iter13_reg <= p_read_56_reg_3224_pp0_iter12_reg;
            p_read_56_reg_3224_pp0_iter14_reg <= p_read_56_reg_3224_pp0_iter13_reg;
            p_read_56_reg_3224_pp0_iter15_reg <= p_read_56_reg_3224_pp0_iter14_reg;
            p_read_56_reg_3224_pp0_iter16_reg <= p_read_56_reg_3224_pp0_iter15_reg;
            p_read_56_reg_3224_pp0_iter17_reg <= p_read_56_reg_3224_pp0_iter16_reg;
            p_read_56_reg_3224_pp0_iter18_reg <= p_read_56_reg_3224_pp0_iter17_reg;
            p_read_56_reg_3224_pp0_iter19_reg <= p_read_56_reg_3224_pp0_iter18_reg;
            p_read_56_reg_3224_pp0_iter1_reg <= p_read_56_reg_3224;
            p_read_56_reg_3224_pp0_iter20_reg <= p_read_56_reg_3224_pp0_iter19_reg;
            p_read_56_reg_3224_pp0_iter21_reg <= p_read_56_reg_3224_pp0_iter20_reg;
            p_read_56_reg_3224_pp0_iter22_reg <= p_read_56_reg_3224_pp0_iter21_reg;
            p_read_56_reg_3224_pp0_iter23_reg <= p_read_56_reg_3224_pp0_iter22_reg;
            p_read_56_reg_3224_pp0_iter24_reg <= p_read_56_reg_3224_pp0_iter23_reg;
            p_read_56_reg_3224_pp0_iter25_reg <= p_read_56_reg_3224_pp0_iter24_reg;
            p_read_56_reg_3224_pp0_iter26_reg <= p_read_56_reg_3224_pp0_iter25_reg;
            p_read_56_reg_3224_pp0_iter27_reg <= p_read_56_reg_3224_pp0_iter26_reg;
            p_read_56_reg_3224_pp0_iter28_reg <= p_read_56_reg_3224_pp0_iter27_reg;
            p_read_56_reg_3224_pp0_iter29_reg <= p_read_56_reg_3224_pp0_iter28_reg;
            p_read_56_reg_3224_pp0_iter2_reg <= p_read_56_reg_3224_pp0_iter1_reg;
            p_read_56_reg_3224_pp0_iter30_reg <= p_read_56_reg_3224_pp0_iter29_reg;
            p_read_56_reg_3224_pp0_iter31_reg <= p_read_56_reg_3224_pp0_iter30_reg;
            p_read_56_reg_3224_pp0_iter32_reg <= p_read_56_reg_3224_pp0_iter31_reg;
            p_read_56_reg_3224_pp0_iter33_reg <= p_read_56_reg_3224_pp0_iter32_reg;
            p_read_56_reg_3224_pp0_iter34_reg <= p_read_56_reg_3224_pp0_iter33_reg;
            p_read_56_reg_3224_pp0_iter35_reg <= p_read_56_reg_3224_pp0_iter34_reg;
            p_read_56_reg_3224_pp0_iter36_reg <= p_read_56_reg_3224_pp0_iter35_reg;
            p_read_56_reg_3224_pp0_iter37_reg <= p_read_56_reg_3224_pp0_iter36_reg;
            p_read_56_reg_3224_pp0_iter38_reg <= p_read_56_reg_3224_pp0_iter37_reg;
            p_read_56_reg_3224_pp0_iter39_reg <= p_read_56_reg_3224_pp0_iter38_reg;
            p_read_56_reg_3224_pp0_iter3_reg <= p_read_56_reg_3224_pp0_iter2_reg;
            p_read_56_reg_3224_pp0_iter40_reg <= p_read_56_reg_3224_pp0_iter39_reg;
            p_read_56_reg_3224_pp0_iter41_reg <= p_read_56_reg_3224_pp0_iter40_reg;
            p_read_56_reg_3224_pp0_iter42_reg <= p_read_56_reg_3224_pp0_iter41_reg;
            p_read_56_reg_3224_pp0_iter43_reg <= p_read_56_reg_3224_pp0_iter42_reg;
            p_read_56_reg_3224_pp0_iter44_reg <= p_read_56_reg_3224_pp0_iter43_reg;
            p_read_56_reg_3224_pp0_iter45_reg <= p_read_56_reg_3224_pp0_iter44_reg;
            p_read_56_reg_3224_pp0_iter46_reg <= p_read_56_reg_3224_pp0_iter45_reg;
            p_read_56_reg_3224_pp0_iter47_reg <= p_read_56_reg_3224_pp0_iter46_reg;
            p_read_56_reg_3224_pp0_iter48_reg <= p_read_56_reg_3224_pp0_iter47_reg;
            p_read_56_reg_3224_pp0_iter49_reg <= p_read_56_reg_3224_pp0_iter48_reg;
            p_read_56_reg_3224_pp0_iter4_reg <= p_read_56_reg_3224_pp0_iter3_reg;
            p_read_56_reg_3224_pp0_iter50_reg <= p_read_56_reg_3224_pp0_iter49_reg;
            p_read_56_reg_3224_pp0_iter51_reg <= p_read_56_reg_3224_pp0_iter50_reg;
            p_read_56_reg_3224_pp0_iter52_reg <= p_read_56_reg_3224_pp0_iter51_reg;
            p_read_56_reg_3224_pp0_iter53_reg <= p_read_56_reg_3224_pp0_iter52_reg;
            p_read_56_reg_3224_pp0_iter54_reg <= p_read_56_reg_3224_pp0_iter53_reg;
            p_read_56_reg_3224_pp0_iter55_reg <= p_read_56_reg_3224_pp0_iter54_reg;
            p_read_56_reg_3224_pp0_iter56_reg <= p_read_56_reg_3224_pp0_iter55_reg;
            p_read_56_reg_3224_pp0_iter57_reg <= p_read_56_reg_3224_pp0_iter56_reg;
            p_read_56_reg_3224_pp0_iter58_reg <= p_read_56_reg_3224_pp0_iter57_reg;
            p_read_56_reg_3224_pp0_iter59_reg <= p_read_56_reg_3224_pp0_iter58_reg;
            p_read_56_reg_3224_pp0_iter5_reg <= p_read_56_reg_3224_pp0_iter4_reg;
            p_read_56_reg_3224_pp0_iter60_reg <= p_read_56_reg_3224_pp0_iter59_reg;
            p_read_56_reg_3224_pp0_iter61_reg <= p_read_56_reg_3224_pp0_iter60_reg;
            p_read_56_reg_3224_pp0_iter62_reg <= p_read_56_reg_3224_pp0_iter61_reg;
            p_read_56_reg_3224_pp0_iter63_reg <= p_read_56_reg_3224_pp0_iter62_reg;
            p_read_56_reg_3224_pp0_iter64_reg <= p_read_56_reg_3224_pp0_iter63_reg;
            p_read_56_reg_3224_pp0_iter65_reg <= p_read_56_reg_3224_pp0_iter64_reg;
            p_read_56_reg_3224_pp0_iter66_reg <= p_read_56_reg_3224_pp0_iter65_reg;
            p_read_56_reg_3224_pp0_iter67_reg <= p_read_56_reg_3224_pp0_iter66_reg;
            p_read_56_reg_3224_pp0_iter68_reg <= p_read_56_reg_3224_pp0_iter67_reg;
            p_read_56_reg_3224_pp0_iter69_reg <= p_read_56_reg_3224_pp0_iter68_reg;
            p_read_56_reg_3224_pp0_iter6_reg <= p_read_56_reg_3224_pp0_iter5_reg;
            p_read_56_reg_3224_pp0_iter70_reg <= p_read_56_reg_3224_pp0_iter69_reg;
            p_read_56_reg_3224_pp0_iter71_reg <= p_read_56_reg_3224_pp0_iter70_reg;
            p_read_56_reg_3224_pp0_iter72_reg <= p_read_56_reg_3224_pp0_iter71_reg;
            p_read_56_reg_3224_pp0_iter73_reg <= p_read_56_reg_3224_pp0_iter72_reg;
            p_read_56_reg_3224_pp0_iter74_reg <= p_read_56_reg_3224_pp0_iter73_reg;
            p_read_56_reg_3224_pp0_iter75_reg <= p_read_56_reg_3224_pp0_iter74_reg;
            p_read_56_reg_3224_pp0_iter76_reg <= p_read_56_reg_3224_pp0_iter75_reg;
            p_read_56_reg_3224_pp0_iter7_reg <= p_read_56_reg_3224_pp0_iter6_reg;
            p_read_56_reg_3224_pp0_iter8_reg <= p_read_56_reg_3224_pp0_iter7_reg;
            p_read_56_reg_3224_pp0_iter9_reg <= p_read_56_reg_3224_pp0_iter8_reg;
            p_read_57_reg_3229 <= p_read7_int_reg;
            p_read_57_reg_3229_pp0_iter10_reg <= p_read_57_reg_3229_pp0_iter9_reg;
            p_read_57_reg_3229_pp0_iter11_reg <= p_read_57_reg_3229_pp0_iter10_reg;
            p_read_57_reg_3229_pp0_iter12_reg <= p_read_57_reg_3229_pp0_iter11_reg;
            p_read_57_reg_3229_pp0_iter13_reg <= p_read_57_reg_3229_pp0_iter12_reg;
            p_read_57_reg_3229_pp0_iter14_reg <= p_read_57_reg_3229_pp0_iter13_reg;
            p_read_57_reg_3229_pp0_iter15_reg <= p_read_57_reg_3229_pp0_iter14_reg;
            p_read_57_reg_3229_pp0_iter16_reg <= p_read_57_reg_3229_pp0_iter15_reg;
            p_read_57_reg_3229_pp0_iter17_reg <= p_read_57_reg_3229_pp0_iter16_reg;
            p_read_57_reg_3229_pp0_iter18_reg <= p_read_57_reg_3229_pp0_iter17_reg;
            p_read_57_reg_3229_pp0_iter19_reg <= p_read_57_reg_3229_pp0_iter18_reg;
            p_read_57_reg_3229_pp0_iter1_reg <= p_read_57_reg_3229;
            p_read_57_reg_3229_pp0_iter20_reg <= p_read_57_reg_3229_pp0_iter19_reg;
            p_read_57_reg_3229_pp0_iter21_reg <= p_read_57_reg_3229_pp0_iter20_reg;
            p_read_57_reg_3229_pp0_iter22_reg <= p_read_57_reg_3229_pp0_iter21_reg;
            p_read_57_reg_3229_pp0_iter23_reg <= p_read_57_reg_3229_pp0_iter22_reg;
            p_read_57_reg_3229_pp0_iter24_reg <= p_read_57_reg_3229_pp0_iter23_reg;
            p_read_57_reg_3229_pp0_iter25_reg <= p_read_57_reg_3229_pp0_iter24_reg;
            p_read_57_reg_3229_pp0_iter26_reg <= p_read_57_reg_3229_pp0_iter25_reg;
            p_read_57_reg_3229_pp0_iter27_reg <= p_read_57_reg_3229_pp0_iter26_reg;
            p_read_57_reg_3229_pp0_iter28_reg <= p_read_57_reg_3229_pp0_iter27_reg;
            p_read_57_reg_3229_pp0_iter29_reg <= p_read_57_reg_3229_pp0_iter28_reg;
            p_read_57_reg_3229_pp0_iter2_reg <= p_read_57_reg_3229_pp0_iter1_reg;
            p_read_57_reg_3229_pp0_iter30_reg <= p_read_57_reg_3229_pp0_iter29_reg;
            p_read_57_reg_3229_pp0_iter31_reg <= p_read_57_reg_3229_pp0_iter30_reg;
            p_read_57_reg_3229_pp0_iter32_reg <= p_read_57_reg_3229_pp0_iter31_reg;
            p_read_57_reg_3229_pp0_iter33_reg <= p_read_57_reg_3229_pp0_iter32_reg;
            p_read_57_reg_3229_pp0_iter34_reg <= p_read_57_reg_3229_pp0_iter33_reg;
            p_read_57_reg_3229_pp0_iter35_reg <= p_read_57_reg_3229_pp0_iter34_reg;
            p_read_57_reg_3229_pp0_iter36_reg <= p_read_57_reg_3229_pp0_iter35_reg;
            p_read_57_reg_3229_pp0_iter37_reg <= p_read_57_reg_3229_pp0_iter36_reg;
            p_read_57_reg_3229_pp0_iter38_reg <= p_read_57_reg_3229_pp0_iter37_reg;
            p_read_57_reg_3229_pp0_iter39_reg <= p_read_57_reg_3229_pp0_iter38_reg;
            p_read_57_reg_3229_pp0_iter3_reg <= p_read_57_reg_3229_pp0_iter2_reg;
            p_read_57_reg_3229_pp0_iter40_reg <= p_read_57_reg_3229_pp0_iter39_reg;
            p_read_57_reg_3229_pp0_iter41_reg <= p_read_57_reg_3229_pp0_iter40_reg;
            p_read_57_reg_3229_pp0_iter42_reg <= p_read_57_reg_3229_pp0_iter41_reg;
            p_read_57_reg_3229_pp0_iter43_reg <= p_read_57_reg_3229_pp0_iter42_reg;
            p_read_57_reg_3229_pp0_iter44_reg <= p_read_57_reg_3229_pp0_iter43_reg;
            p_read_57_reg_3229_pp0_iter45_reg <= p_read_57_reg_3229_pp0_iter44_reg;
            p_read_57_reg_3229_pp0_iter46_reg <= p_read_57_reg_3229_pp0_iter45_reg;
            p_read_57_reg_3229_pp0_iter47_reg <= p_read_57_reg_3229_pp0_iter46_reg;
            p_read_57_reg_3229_pp0_iter48_reg <= p_read_57_reg_3229_pp0_iter47_reg;
            p_read_57_reg_3229_pp0_iter49_reg <= p_read_57_reg_3229_pp0_iter48_reg;
            p_read_57_reg_3229_pp0_iter4_reg <= p_read_57_reg_3229_pp0_iter3_reg;
            p_read_57_reg_3229_pp0_iter50_reg <= p_read_57_reg_3229_pp0_iter49_reg;
            p_read_57_reg_3229_pp0_iter51_reg <= p_read_57_reg_3229_pp0_iter50_reg;
            p_read_57_reg_3229_pp0_iter52_reg <= p_read_57_reg_3229_pp0_iter51_reg;
            p_read_57_reg_3229_pp0_iter53_reg <= p_read_57_reg_3229_pp0_iter52_reg;
            p_read_57_reg_3229_pp0_iter54_reg <= p_read_57_reg_3229_pp0_iter53_reg;
            p_read_57_reg_3229_pp0_iter55_reg <= p_read_57_reg_3229_pp0_iter54_reg;
            p_read_57_reg_3229_pp0_iter56_reg <= p_read_57_reg_3229_pp0_iter55_reg;
            p_read_57_reg_3229_pp0_iter57_reg <= p_read_57_reg_3229_pp0_iter56_reg;
            p_read_57_reg_3229_pp0_iter58_reg <= p_read_57_reg_3229_pp0_iter57_reg;
            p_read_57_reg_3229_pp0_iter59_reg <= p_read_57_reg_3229_pp0_iter58_reg;
            p_read_57_reg_3229_pp0_iter5_reg <= p_read_57_reg_3229_pp0_iter4_reg;
            p_read_57_reg_3229_pp0_iter60_reg <= p_read_57_reg_3229_pp0_iter59_reg;
            p_read_57_reg_3229_pp0_iter61_reg <= p_read_57_reg_3229_pp0_iter60_reg;
            p_read_57_reg_3229_pp0_iter62_reg <= p_read_57_reg_3229_pp0_iter61_reg;
            p_read_57_reg_3229_pp0_iter63_reg <= p_read_57_reg_3229_pp0_iter62_reg;
            p_read_57_reg_3229_pp0_iter64_reg <= p_read_57_reg_3229_pp0_iter63_reg;
            p_read_57_reg_3229_pp0_iter65_reg <= p_read_57_reg_3229_pp0_iter64_reg;
            p_read_57_reg_3229_pp0_iter66_reg <= p_read_57_reg_3229_pp0_iter65_reg;
            p_read_57_reg_3229_pp0_iter67_reg <= p_read_57_reg_3229_pp0_iter66_reg;
            p_read_57_reg_3229_pp0_iter68_reg <= p_read_57_reg_3229_pp0_iter67_reg;
            p_read_57_reg_3229_pp0_iter69_reg <= p_read_57_reg_3229_pp0_iter68_reg;
            p_read_57_reg_3229_pp0_iter6_reg <= p_read_57_reg_3229_pp0_iter5_reg;
            p_read_57_reg_3229_pp0_iter70_reg <= p_read_57_reg_3229_pp0_iter69_reg;
            p_read_57_reg_3229_pp0_iter71_reg <= p_read_57_reg_3229_pp0_iter70_reg;
            p_read_57_reg_3229_pp0_iter72_reg <= p_read_57_reg_3229_pp0_iter71_reg;
            p_read_57_reg_3229_pp0_iter73_reg <= p_read_57_reg_3229_pp0_iter72_reg;
            p_read_57_reg_3229_pp0_iter74_reg <= p_read_57_reg_3229_pp0_iter73_reg;
            p_read_57_reg_3229_pp0_iter75_reg <= p_read_57_reg_3229_pp0_iter74_reg;
            p_read_57_reg_3229_pp0_iter76_reg <= p_read_57_reg_3229_pp0_iter75_reg;
            p_read_57_reg_3229_pp0_iter7_reg <= p_read_57_reg_3229_pp0_iter6_reg;
            p_read_57_reg_3229_pp0_iter8_reg <= p_read_57_reg_3229_pp0_iter7_reg;
            p_read_57_reg_3229_pp0_iter9_reg <= p_read_57_reg_3229_pp0_iter8_reg;
            p_read_58_reg_3234 <= p_read6_int_reg;
            p_read_58_reg_3234_pp0_iter10_reg <= p_read_58_reg_3234_pp0_iter9_reg;
            p_read_58_reg_3234_pp0_iter11_reg <= p_read_58_reg_3234_pp0_iter10_reg;
            p_read_58_reg_3234_pp0_iter12_reg <= p_read_58_reg_3234_pp0_iter11_reg;
            p_read_58_reg_3234_pp0_iter13_reg <= p_read_58_reg_3234_pp0_iter12_reg;
            p_read_58_reg_3234_pp0_iter14_reg <= p_read_58_reg_3234_pp0_iter13_reg;
            p_read_58_reg_3234_pp0_iter15_reg <= p_read_58_reg_3234_pp0_iter14_reg;
            p_read_58_reg_3234_pp0_iter16_reg <= p_read_58_reg_3234_pp0_iter15_reg;
            p_read_58_reg_3234_pp0_iter17_reg <= p_read_58_reg_3234_pp0_iter16_reg;
            p_read_58_reg_3234_pp0_iter18_reg <= p_read_58_reg_3234_pp0_iter17_reg;
            p_read_58_reg_3234_pp0_iter19_reg <= p_read_58_reg_3234_pp0_iter18_reg;
            p_read_58_reg_3234_pp0_iter1_reg <= p_read_58_reg_3234;
            p_read_58_reg_3234_pp0_iter20_reg <= p_read_58_reg_3234_pp0_iter19_reg;
            p_read_58_reg_3234_pp0_iter21_reg <= p_read_58_reg_3234_pp0_iter20_reg;
            p_read_58_reg_3234_pp0_iter22_reg <= p_read_58_reg_3234_pp0_iter21_reg;
            p_read_58_reg_3234_pp0_iter23_reg <= p_read_58_reg_3234_pp0_iter22_reg;
            p_read_58_reg_3234_pp0_iter24_reg <= p_read_58_reg_3234_pp0_iter23_reg;
            p_read_58_reg_3234_pp0_iter25_reg <= p_read_58_reg_3234_pp0_iter24_reg;
            p_read_58_reg_3234_pp0_iter26_reg <= p_read_58_reg_3234_pp0_iter25_reg;
            p_read_58_reg_3234_pp0_iter27_reg <= p_read_58_reg_3234_pp0_iter26_reg;
            p_read_58_reg_3234_pp0_iter28_reg <= p_read_58_reg_3234_pp0_iter27_reg;
            p_read_58_reg_3234_pp0_iter29_reg <= p_read_58_reg_3234_pp0_iter28_reg;
            p_read_58_reg_3234_pp0_iter2_reg <= p_read_58_reg_3234_pp0_iter1_reg;
            p_read_58_reg_3234_pp0_iter30_reg <= p_read_58_reg_3234_pp0_iter29_reg;
            p_read_58_reg_3234_pp0_iter31_reg <= p_read_58_reg_3234_pp0_iter30_reg;
            p_read_58_reg_3234_pp0_iter32_reg <= p_read_58_reg_3234_pp0_iter31_reg;
            p_read_58_reg_3234_pp0_iter33_reg <= p_read_58_reg_3234_pp0_iter32_reg;
            p_read_58_reg_3234_pp0_iter34_reg <= p_read_58_reg_3234_pp0_iter33_reg;
            p_read_58_reg_3234_pp0_iter35_reg <= p_read_58_reg_3234_pp0_iter34_reg;
            p_read_58_reg_3234_pp0_iter36_reg <= p_read_58_reg_3234_pp0_iter35_reg;
            p_read_58_reg_3234_pp0_iter37_reg <= p_read_58_reg_3234_pp0_iter36_reg;
            p_read_58_reg_3234_pp0_iter38_reg <= p_read_58_reg_3234_pp0_iter37_reg;
            p_read_58_reg_3234_pp0_iter39_reg <= p_read_58_reg_3234_pp0_iter38_reg;
            p_read_58_reg_3234_pp0_iter3_reg <= p_read_58_reg_3234_pp0_iter2_reg;
            p_read_58_reg_3234_pp0_iter40_reg <= p_read_58_reg_3234_pp0_iter39_reg;
            p_read_58_reg_3234_pp0_iter41_reg <= p_read_58_reg_3234_pp0_iter40_reg;
            p_read_58_reg_3234_pp0_iter42_reg <= p_read_58_reg_3234_pp0_iter41_reg;
            p_read_58_reg_3234_pp0_iter43_reg <= p_read_58_reg_3234_pp0_iter42_reg;
            p_read_58_reg_3234_pp0_iter44_reg <= p_read_58_reg_3234_pp0_iter43_reg;
            p_read_58_reg_3234_pp0_iter45_reg <= p_read_58_reg_3234_pp0_iter44_reg;
            p_read_58_reg_3234_pp0_iter46_reg <= p_read_58_reg_3234_pp0_iter45_reg;
            p_read_58_reg_3234_pp0_iter47_reg <= p_read_58_reg_3234_pp0_iter46_reg;
            p_read_58_reg_3234_pp0_iter48_reg <= p_read_58_reg_3234_pp0_iter47_reg;
            p_read_58_reg_3234_pp0_iter49_reg <= p_read_58_reg_3234_pp0_iter48_reg;
            p_read_58_reg_3234_pp0_iter4_reg <= p_read_58_reg_3234_pp0_iter3_reg;
            p_read_58_reg_3234_pp0_iter50_reg <= p_read_58_reg_3234_pp0_iter49_reg;
            p_read_58_reg_3234_pp0_iter51_reg <= p_read_58_reg_3234_pp0_iter50_reg;
            p_read_58_reg_3234_pp0_iter52_reg <= p_read_58_reg_3234_pp0_iter51_reg;
            p_read_58_reg_3234_pp0_iter53_reg <= p_read_58_reg_3234_pp0_iter52_reg;
            p_read_58_reg_3234_pp0_iter54_reg <= p_read_58_reg_3234_pp0_iter53_reg;
            p_read_58_reg_3234_pp0_iter55_reg <= p_read_58_reg_3234_pp0_iter54_reg;
            p_read_58_reg_3234_pp0_iter56_reg <= p_read_58_reg_3234_pp0_iter55_reg;
            p_read_58_reg_3234_pp0_iter57_reg <= p_read_58_reg_3234_pp0_iter56_reg;
            p_read_58_reg_3234_pp0_iter58_reg <= p_read_58_reg_3234_pp0_iter57_reg;
            p_read_58_reg_3234_pp0_iter59_reg <= p_read_58_reg_3234_pp0_iter58_reg;
            p_read_58_reg_3234_pp0_iter5_reg <= p_read_58_reg_3234_pp0_iter4_reg;
            p_read_58_reg_3234_pp0_iter60_reg <= p_read_58_reg_3234_pp0_iter59_reg;
            p_read_58_reg_3234_pp0_iter61_reg <= p_read_58_reg_3234_pp0_iter60_reg;
            p_read_58_reg_3234_pp0_iter62_reg <= p_read_58_reg_3234_pp0_iter61_reg;
            p_read_58_reg_3234_pp0_iter63_reg <= p_read_58_reg_3234_pp0_iter62_reg;
            p_read_58_reg_3234_pp0_iter64_reg <= p_read_58_reg_3234_pp0_iter63_reg;
            p_read_58_reg_3234_pp0_iter65_reg <= p_read_58_reg_3234_pp0_iter64_reg;
            p_read_58_reg_3234_pp0_iter66_reg <= p_read_58_reg_3234_pp0_iter65_reg;
            p_read_58_reg_3234_pp0_iter67_reg <= p_read_58_reg_3234_pp0_iter66_reg;
            p_read_58_reg_3234_pp0_iter68_reg <= p_read_58_reg_3234_pp0_iter67_reg;
            p_read_58_reg_3234_pp0_iter69_reg <= p_read_58_reg_3234_pp0_iter68_reg;
            p_read_58_reg_3234_pp0_iter6_reg <= p_read_58_reg_3234_pp0_iter5_reg;
            p_read_58_reg_3234_pp0_iter70_reg <= p_read_58_reg_3234_pp0_iter69_reg;
            p_read_58_reg_3234_pp0_iter71_reg <= p_read_58_reg_3234_pp0_iter70_reg;
            p_read_58_reg_3234_pp0_iter72_reg <= p_read_58_reg_3234_pp0_iter71_reg;
            p_read_58_reg_3234_pp0_iter73_reg <= p_read_58_reg_3234_pp0_iter72_reg;
            p_read_58_reg_3234_pp0_iter74_reg <= p_read_58_reg_3234_pp0_iter73_reg;
            p_read_58_reg_3234_pp0_iter75_reg <= p_read_58_reg_3234_pp0_iter74_reg;
            p_read_58_reg_3234_pp0_iter76_reg <= p_read_58_reg_3234_pp0_iter75_reg;
            p_read_58_reg_3234_pp0_iter7_reg <= p_read_58_reg_3234_pp0_iter6_reg;
            p_read_58_reg_3234_pp0_iter8_reg <= p_read_58_reg_3234_pp0_iter7_reg;
            p_read_58_reg_3234_pp0_iter9_reg <= p_read_58_reg_3234_pp0_iter8_reg;
            p_read_59_reg_3239 <= p_read5_int_reg;
            p_read_59_reg_3239_pp0_iter10_reg <= p_read_59_reg_3239_pp0_iter9_reg;
            p_read_59_reg_3239_pp0_iter11_reg <= p_read_59_reg_3239_pp0_iter10_reg;
            p_read_59_reg_3239_pp0_iter12_reg <= p_read_59_reg_3239_pp0_iter11_reg;
            p_read_59_reg_3239_pp0_iter13_reg <= p_read_59_reg_3239_pp0_iter12_reg;
            p_read_59_reg_3239_pp0_iter14_reg <= p_read_59_reg_3239_pp0_iter13_reg;
            p_read_59_reg_3239_pp0_iter15_reg <= p_read_59_reg_3239_pp0_iter14_reg;
            p_read_59_reg_3239_pp0_iter16_reg <= p_read_59_reg_3239_pp0_iter15_reg;
            p_read_59_reg_3239_pp0_iter17_reg <= p_read_59_reg_3239_pp0_iter16_reg;
            p_read_59_reg_3239_pp0_iter18_reg <= p_read_59_reg_3239_pp0_iter17_reg;
            p_read_59_reg_3239_pp0_iter19_reg <= p_read_59_reg_3239_pp0_iter18_reg;
            p_read_59_reg_3239_pp0_iter1_reg <= p_read_59_reg_3239;
            p_read_59_reg_3239_pp0_iter20_reg <= p_read_59_reg_3239_pp0_iter19_reg;
            p_read_59_reg_3239_pp0_iter21_reg <= p_read_59_reg_3239_pp0_iter20_reg;
            p_read_59_reg_3239_pp0_iter22_reg <= p_read_59_reg_3239_pp0_iter21_reg;
            p_read_59_reg_3239_pp0_iter23_reg <= p_read_59_reg_3239_pp0_iter22_reg;
            p_read_59_reg_3239_pp0_iter24_reg <= p_read_59_reg_3239_pp0_iter23_reg;
            p_read_59_reg_3239_pp0_iter25_reg <= p_read_59_reg_3239_pp0_iter24_reg;
            p_read_59_reg_3239_pp0_iter26_reg <= p_read_59_reg_3239_pp0_iter25_reg;
            p_read_59_reg_3239_pp0_iter27_reg <= p_read_59_reg_3239_pp0_iter26_reg;
            p_read_59_reg_3239_pp0_iter28_reg <= p_read_59_reg_3239_pp0_iter27_reg;
            p_read_59_reg_3239_pp0_iter29_reg <= p_read_59_reg_3239_pp0_iter28_reg;
            p_read_59_reg_3239_pp0_iter2_reg <= p_read_59_reg_3239_pp0_iter1_reg;
            p_read_59_reg_3239_pp0_iter30_reg <= p_read_59_reg_3239_pp0_iter29_reg;
            p_read_59_reg_3239_pp0_iter31_reg <= p_read_59_reg_3239_pp0_iter30_reg;
            p_read_59_reg_3239_pp0_iter32_reg <= p_read_59_reg_3239_pp0_iter31_reg;
            p_read_59_reg_3239_pp0_iter33_reg <= p_read_59_reg_3239_pp0_iter32_reg;
            p_read_59_reg_3239_pp0_iter34_reg <= p_read_59_reg_3239_pp0_iter33_reg;
            p_read_59_reg_3239_pp0_iter35_reg <= p_read_59_reg_3239_pp0_iter34_reg;
            p_read_59_reg_3239_pp0_iter36_reg <= p_read_59_reg_3239_pp0_iter35_reg;
            p_read_59_reg_3239_pp0_iter37_reg <= p_read_59_reg_3239_pp0_iter36_reg;
            p_read_59_reg_3239_pp0_iter38_reg <= p_read_59_reg_3239_pp0_iter37_reg;
            p_read_59_reg_3239_pp0_iter39_reg <= p_read_59_reg_3239_pp0_iter38_reg;
            p_read_59_reg_3239_pp0_iter3_reg <= p_read_59_reg_3239_pp0_iter2_reg;
            p_read_59_reg_3239_pp0_iter40_reg <= p_read_59_reg_3239_pp0_iter39_reg;
            p_read_59_reg_3239_pp0_iter41_reg <= p_read_59_reg_3239_pp0_iter40_reg;
            p_read_59_reg_3239_pp0_iter42_reg <= p_read_59_reg_3239_pp0_iter41_reg;
            p_read_59_reg_3239_pp0_iter43_reg <= p_read_59_reg_3239_pp0_iter42_reg;
            p_read_59_reg_3239_pp0_iter44_reg <= p_read_59_reg_3239_pp0_iter43_reg;
            p_read_59_reg_3239_pp0_iter45_reg <= p_read_59_reg_3239_pp0_iter44_reg;
            p_read_59_reg_3239_pp0_iter46_reg <= p_read_59_reg_3239_pp0_iter45_reg;
            p_read_59_reg_3239_pp0_iter47_reg <= p_read_59_reg_3239_pp0_iter46_reg;
            p_read_59_reg_3239_pp0_iter48_reg <= p_read_59_reg_3239_pp0_iter47_reg;
            p_read_59_reg_3239_pp0_iter49_reg <= p_read_59_reg_3239_pp0_iter48_reg;
            p_read_59_reg_3239_pp0_iter4_reg <= p_read_59_reg_3239_pp0_iter3_reg;
            p_read_59_reg_3239_pp0_iter50_reg <= p_read_59_reg_3239_pp0_iter49_reg;
            p_read_59_reg_3239_pp0_iter51_reg <= p_read_59_reg_3239_pp0_iter50_reg;
            p_read_59_reg_3239_pp0_iter52_reg <= p_read_59_reg_3239_pp0_iter51_reg;
            p_read_59_reg_3239_pp0_iter53_reg <= p_read_59_reg_3239_pp0_iter52_reg;
            p_read_59_reg_3239_pp0_iter54_reg <= p_read_59_reg_3239_pp0_iter53_reg;
            p_read_59_reg_3239_pp0_iter55_reg <= p_read_59_reg_3239_pp0_iter54_reg;
            p_read_59_reg_3239_pp0_iter56_reg <= p_read_59_reg_3239_pp0_iter55_reg;
            p_read_59_reg_3239_pp0_iter57_reg <= p_read_59_reg_3239_pp0_iter56_reg;
            p_read_59_reg_3239_pp0_iter58_reg <= p_read_59_reg_3239_pp0_iter57_reg;
            p_read_59_reg_3239_pp0_iter59_reg <= p_read_59_reg_3239_pp0_iter58_reg;
            p_read_59_reg_3239_pp0_iter5_reg <= p_read_59_reg_3239_pp0_iter4_reg;
            p_read_59_reg_3239_pp0_iter60_reg <= p_read_59_reg_3239_pp0_iter59_reg;
            p_read_59_reg_3239_pp0_iter61_reg <= p_read_59_reg_3239_pp0_iter60_reg;
            p_read_59_reg_3239_pp0_iter62_reg <= p_read_59_reg_3239_pp0_iter61_reg;
            p_read_59_reg_3239_pp0_iter63_reg <= p_read_59_reg_3239_pp0_iter62_reg;
            p_read_59_reg_3239_pp0_iter64_reg <= p_read_59_reg_3239_pp0_iter63_reg;
            p_read_59_reg_3239_pp0_iter65_reg <= p_read_59_reg_3239_pp0_iter64_reg;
            p_read_59_reg_3239_pp0_iter66_reg <= p_read_59_reg_3239_pp0_iter65_reg;
            p_read_59_reg_3239_pp0_iter67_reg <= p_read_59_reg_3239_pp0_iter66_reg;
            p_read_59_reg_3239_pp0_iter68_reg <= p_read_59_reg_3239_pp0_iter67_reg;
            p_read_59_reg_3239_pp0_iter69_reg <= p_read_59_reg_3239_pp0_iter68_reg;
            p_read_59_reg_3239_pp0_iter6_reg <= p_read_59_reg_3239_pp0_iter5_reg;
            p_read_59_reg_3239_pp0_iter70_reg <= p_read_59_reg_3239_pp0_iter69_reg;
            p_read_59_reg_3239_pp0_iter71_reg <= p_read_59_reg_3239_pp0_iter70_reg;
            p_read_59_reg_3239_pp0_iter72_reg <= p_read_59_reg_3239_pp0_iter71_reg;
            p_read_59_reg_3239_pp0_iter73_reg <= p_read_59_reg_3239_pp0_iter72_reg;
            p_read_59_reg_3239_pp0_iter74_reg <= p_read_59_reg_3239_pp0_iter73_reg;
            p_read_59_reg_3239_pp0_iter75_reg <= p_read_59_reg_3239_pp0_iter74_reg;
            p_read_59_reg_3239_pp0_iter76_reg <= p_read_59_reg_3239_pp0_iter75_reg;
            p_read_59_reg_3239_pp0_iter7_reg <= p_read_59_reg_3239_pp0_iter6_reg;
            p_read_59_reg_3239_pp0_iter8_reg <= p_read_59_reg_3239_pp0_iter7_reg;
            p_read_59_reg_3239_pp0_iter9_reg <= p_read_59_reg_3239_pp0_iter8_reg;
            p_read_60_reg_3244 <= p_read4_int_reg;
            p_read_60_reg_3244_pp0_iter10_reg <= p_read_60_reg_3244_pp0_iter9_reg;
            p_read_60_reg_3244_pp0_iter11_reg <= p_read_60_reg_3244_pp0_iter10_reg;
            p_read_60_reg_3244_pp0_iter12_reg <= p_read_60_reg_3244_pp0_iter11_reg;
            p_read_60_reg_3244_pp0_iter13_reg <= p_read_60_reg_3244_pp0_iter12_reg;
            p_read_60_reg_3244_pp0_iter14_reg <= p_read_60_reg_3244_pp0_iter13_reg;
            p_read_60_reg_3244_pp0_iter15_reg <= p_read_60_reg_3244_pp0_iter14_reg;
            p_read_60_reg_3244_pp0_iter16_reg <= p_read_60_reg_3244_pp0_iter15_reg;
            p_read_60_reg_3244_pp0_iter17_reg <= p_read_60_reg_3244_pp0_iter16_reg;
            p_read_60_reg_3244_pp0_iter18_reg <= p_read_60_reg_3244_pp0_iter17_reg;
            p_read_60_reg_3244_pp0_iter19_reg <= p_read_60_reg_3244_pp0_iter18_reg;
            p_read_60_reg_3244_pp0_iter1_reg <= p_read_60_reg_3244;
            p_read_60_reg_3244_pp0_iter20_reg <= p_read_60_reg_3244_pp0_iter19_reg;
            p_read_60_reg_3244_pp0_iter21_reg <= p_read_60_reg_3244_pp0_iter20_reg;
            p_read_60_reg_3244_pp0_iter22_reg <= p_read_60_reg_3244_pp0_iter21_reg;
            p_read_60_reg_3244_pp0_iter23_reg <= p_read_60_reg_3244_pp0_iter22_reg;
            p_read_60_reg_3244_pp0_iter24_reg <= p_read_60_reg_3244_pp0_iter23_reg;
            p_read_60_reg_3244_pp0_iter25_reg <= p_read_60_reg_3244_pp0_iter24_reg;
            p_read_60_reg_3244_pp0_iter26_reg <= p_read_60_reg_3244_pp0_iter25_reg;
            p_read_60_reg_3244_pp0_iter27_reg <= p_read_60_reg_3244_pp0_iter26_reg;
            p_read_60_reg_3244_pp0_iter28_reg <= p_read_60_reg_3244_pp0_iter27_reg;
            p_read_60_reg_3244_pp0_iter29_reg <= p_read_60_reg_3244_pp0_iter28_reg;
            p_read_60_reg_3244_pp0_iter2_reg <= p_read_60_reg_3244_pp0_iter1_reg;
            p_read_60_reg_3244_pp0_iter30_reg <= p_read_60_reg_3244_pp0_iter29_reg;
            p_read_60_reg_3244_pp0_iter31_reg <= p_read_60_reg_3244_pp0_iter30_reg;
            p_read_60_reg_3244_pp0_iter32_reg <= p_read_60_reg_3244_pp0_iter31_reg;
            p_read_60_reg_3244_pp0_iter33_reg <= p_read_60_reg_3244_pp0_iter32_reg;
            p_read_60_reg_3244_pp0_iter34_reg <= p_read_60_reg_3244_pp0_iter33_reg;
            p_read_60_reg_3244_pp0_iter35_reg <= p_read_60_reg_3244_pp0_iter34_reg;
            p_read_60_reg_3244_pp0_iter36_reg <= p_read_60_reg_3244_pp0_iter35_reg;
            p_read_60_reg_3244_pp0_iter37_reg <= p_read_60_reg_3244_pp0_iter36_reg;
            p_read_60_reg_3244_pp0_iter38_reg <= p_read_60_reg_3244_pp0_iter37_reg;
            p_read_60_reg_3244_pp0_iter39_reg <= p_read_60_reg_3244_pp0_iter38_reg;
            p_read_60_reg_3244_pp0_iter3_reg <= p_read_60_reg_3244_pp0_iter2_reg;
            p_read_60_reg_3244_pp0_iter40_reg <= p_read_60_reg_3244_pp0_iter39_reg;
            p_read_60_reg_3244_pp0_iter41_reg <= p_read_60_reg_3244_pp0_iter40_reg;
            p_read_60_reg_3244_pp0_iter42_reg <= p_read_60_reg_3244_pp0_iter41_reg;
            p_read_60_reg_3244_pp0_iter43_reg <= p_read_60_reg_3244_pp0_iter42_reg;
            p_read_60_reg_3244_pp0_iter44_reg <= p_read_60_reg_3244_pp0_iter43_reg;
            p_read_60_reg_3244_pp0_iter45_reg <= p_read_60_reg_3244_pp0_iter44_reg;
            p_read_60_reg_3244_pp0_iter46_reg <= p_read_60_reg_3244_pp0_iter45_reg;
            p_read_60_reg_3244_pp0_iter47_reg <= p_read_60_reg_3244_pp0_iter46_reg;
            p_read_60_reg_3244_pp0_iter48_reg <= p_read_60_reg_3244_pp0_iter47_reg;
            p_read_60_reg_3244_pp0_iter49_reg <= p_read_60_reg_3244_pp0_iter48_reg;
            p_read_60_reg_3244_pp0_iter4_reg <= p_read_60_reg_3244_pp0_iter3_reg;
            p_read_60_reg_3244_pp0_iter50_reg <= p_read_60_reg_3244_pp0_iter49_reg;
            p_read_60_reg_3244_pp0_iter51_reg <= p_read_60_reg_3244_pp0_iter50_reg;
            p_read_60_reg_3244_pp0_iter52_reg <= p_read_60_reg_3244_pp0_iter51_reg;
            p_read_60_reg_3244_pp0_iter53_reg <= p_read_60_reg_3244_pp0_iter52_reg;
            p_read_60_reg_3244_pp0_iter54_reg <= p_read_60_reg_3244_pp0_iter53_reg;
            p_read_60_reg_3244_pp0_iter55_reg <= p_read_60_reg_3244_pp0_iter54_reg;
            p_read_60_reg_3244_pp0_iter56_reg <= p_read_60_reg_3244_pp0_iter55_reg;
            p_read_60_reg_3244_pp0_iter57_reg <= p_read_60_reg_3244_pp0_iter56_reg;
            p_read_60_reg_3244_pp0_iter58_reg <= p_read_60_reg_3244_pp0_iter57_reg;
            p_read_60_reg_3244_pp0_iter59_reg <= p_read_60_reg_3244_pp0_iter58_reg;
            p_read_60_reg_3244_pp0_iter5_reg <= p_read_60_reg_3244_pp0_iter4_reg;
            p_read_60_reg_3244_pp0_iter60_reg <= p_read_60_reg_3244_pp0_iter59_reg;
            p_read_60_reg_3244_pp0_iter61_reg <= p_read_60_reg_3244_pp0_iter60_reg;
            p_read_60_reg_3244_pp0_iter62_reg <= p_read_60_reg_3244_pp0_iter61_reg;
            p_read_60_reg_3244_pp0_iter63_reg <= p_read_60_reg_3244_pp0_iter62_reg;
            p_read_60_reg_3244_pp0_iter64_reg <= p_read_60_reg_3244_pp0_iter63_reg;
            p_read_60_reg_3244_pp0_iter65_reg <= p_read_60_reg_3244_pp0_iter64_reg;
            p_read_60_reg_3244_pp0_iter66_reg <= p_read_60_reg_3244_pp0_iter65_reg;
            p_read_60_reg_3244_pp0_iter67_reg <= p_read_60_reg_3244_pp0_iter66_reg;
            p_read_60_reg_3244_pp0_iter68_reg <= p_read_60_reg_3244_pp0_iter67_reg;
            p_read_60_reg_3244_pp0_iter69_reg <= p_read_60_reg_3244_pp0_iter68_reg;
            p_read_60_reg_3244_pp0_iter6_reg <= p_read_60_reg_3244_pp0_iter5_reg;
            p_read_60_reg_3244_pp0_iter70_reg <= p_read_60_reg_3244_pp0_iter69_reg;
            p_read_60_reg_3244_pp0_iter71_reg <= p_read_60_reg_3244_pp0_iter70_reg;
            p_read_60_reg_3244_pp0_iter72_reg <= p_read_60_reg_3244_pp0_iter71_reg;
            p_read_60_reg_3244_pp0_iter73_reg <= p_read_60_reg_3244_pp0_iter72_reg;
            p_read_60_reg_3244_pp0_iter74_reg <= p_read_60_reg_3244_pp0_iter73_reg;
            p_read_60_reg_3244_pp0_iter75_reg <= p_read_60_reg_3244_pp0_iter74_reg;
            p_read_60_reg_3244_pp0_iter76_reg <= p_read_60_reg_3244_pp0_iter75_reg;
            p_read_60_reg_3244_pp0_iter7_reg <= p_read_60_reg_3244_pp0_iter6_reg;
            p_read_60_reg_3244_pp0_iter8_reg <= p_read_60_reg_3244_pp0_iter7_reg;
            p_read_60_reg_3244_pp0_iter9_reg <= p_read_60_reg_3244_pp0_iter8_reg;
            p_read_61_reg_3249 <= p_read3_int_reg;
            p_read_61_reg_3249_pp0_iter10_reg <= p_read_61_reg_3249_pp0_iter9_reg;
            p_read_61_reg_3249_pp0_iter11_reg <= p_read_61_reg_3249_pp0_iter10_reg;
            p_read_61_reg_3249_pp0_iter12_reg <= p_read_61_reg_3249_pp0_iter11_reg;
            p_read_61_reg_3249_pp0_iter13_reg <= p_read_61_reg_3249_pp0_iter12_reg;
            p_read_61_reg_3249_pp0_iter14_reg <= p_read_61_reg_3249_pp0_iter13_reg;
            p_read_61_reg_3249_pp0_iter15_reg <= p_read_61_reg_3249_pp0_iter14_reg;
            p_read_61_reg_3249_pp0_iter16_reg <= p_read_61_reg_3249_pp0_iter15_reg;
            p_read_61_reg_3249_pp0_iter17_reg <= p_read_61_reg_3249_pp0_iter16_reg;
            p_read_61_reg_3249_pp0_iter18_reg <= p_read_61_reg_3249_pp0_iter17_reg;
            p_read_61_reg_3249_pp0_iter19_reg <= p_read_61_reg_3249_pp0_iter18_reg;
            p_read_61_reg_3249_pp0_iter1_reg <= p_read_61_reg_3249;
            p_read_61_reg_3249_pp0_iter20_reg <= p_read_61_reg_3249_pp0_iter19_reg;
            p_read_61_reg_3249_pp0_iter21_reg <= p_read_61_reg_3249_pp0_iter20_reg;
            p_read_61_reg_3249_pp0_iter22_reg <= p_read_61_reg_3249_pp0_iter21_reg;
            p_read_61_reg_3249_pp0_iter23_reg <= p_read_61_reg_3249_pp0_iter22_reg;
            p_read_61_reg_3249_pp0_iter24_reg <= p_read_61_reg_3249_pp0_iter23_reg;
            p_read_61_reg_3249_pp0_iter25_reg <= p_read_61_reg_3249_pp0_iter24_reg;
            p_read_61_reg_3249_pp0_iter26_reg <= p_read_61_reg_3249_pp0_iter25_reg;
            p_read_61_reg_3249_pp0_iter27_reg <= p_read_61_reg_3249_pp0_iter26_reg;
            p_read_61_reg_3249_pp0_iter28_reg <= p_read_61_reg_3249_pp0_iter27_reg;
            p_read_61_reg_3249_pp0_iter29_reg <= p_read_61_reg_3249_pp0_iter28_reg;
            p_read_61_reg_3249_pp0_iter2_reg <= p_read_61_reg_3249_pp0_iter1_reg;
            p_read_61_reg_3249_pp0_iter30_reg <= p_read_61_reg_3249_pp0_iter29_reg;
            p_read_61_reg_3249_pp0_iter31_reg <= p_read_61_reg_3249_pp0_iter30_reg;
            p_read_61_reg_3249_pp0_iter32_reg <= p_read_61_reg_3249_pp0_iter31_reg;
            p_read_61_reg_3249_pp0_iter33_reg <= p_read_61_reg_3249_pp0_iter32_reg;
            p_read_61_reg_3249_pp0_iter34_reg <= p_read_61_reg_3249_pp0_iter33_reg;
            p_read_61_reg_3249_pp0_iter35_reg <= p_read_61_reg_3249_pp0_iter34_reg;
            p_read_61_reg_3249_pp0_iter36_reg <= p_read_61_reg_3249_pp0_iter35_reg;
            p_read_61_reg_3249_pp0_iter37_reg <= p_read_61_reg_3249_pp0_iter36_reg;
            p_read_61_reg_3249_pp0_iter38_reg <= p_read_61_reg_3249_pp0_iter37_reg;
            p_read_61_reg_3249_pp0_iter39_reg <= p_read_61_reg_3249_pp0_iter38_reg;
            p_read_61_reg_3249_pp0_iter3_reg <= p_read_61_reg_3249_pp0_iter2_reg;
            p_read_61_reg_3249_pp0_iter40_reg <= p_read_61_reg_3249_pp0_iter39_reg;
            p_read_61_reg_3249_pp0_iter41_reg <= p_read_61_reg_3249_pp0_iter40_reg;
            p_read_61_reg_3249_pp0_iter42_reg <= p_read_61_reg_3249_pp0_iter41_reg;
            p_read_61_reg_3249_pp0_iter43_reg <= p_read_61_reg_3249_pp0_iter42_reg;
            p_read_61_reg_3249_pp0_iter44_reg <= p_read_61_reg_3249_pp0_iter43_reg;
            p_read_61_reg_3249_pp0_iter45_reg <= p_read_61_reg_3249_pp0_iter44_reg;
            p_read_61_reg_3249_pp0_iter46_reg <= p_read_61_reg_3249_pp0_iter45_reg;
            p_read_61_reg_3249_pp0_iter47_reg <= p_read_61_reg_3249_pp0_iter46_reg;
            p_read_61_reg_3249_pp0_iter48_reg <= p_read_61_reg_3249_pp0_iter47_reg;
            p_read_61_reg_3249_pp0_iter49_reg <= p_read_61_reg_3249_pp0_iter48_reg;
            p_read_61_reg_3249_pp0_iter4_reg <= p_read_61_reg_3249_pp0_iter3_reg;
            p_read_61_reg_3249_pp0_iter50_reg <= p_read_61_reg_3249_pp0_iter49_reg;
            p_read_61_reg_3249_pp0_iter51_reg <= p_read_61_reg_3249_pp0_iter50_reg;
            p_read_61_reg_3249_pp0_iter52_reg <= p_read_61_reg_3249_pp0_iter51_reg;
            p_read_61_reg_3249_pp0_iter53_reg <= p_read_61_reg_3249_pp0_iter52_reg;
            p_read_61_reg_3249_pp0_iter54_reg <= p_read_61_reg_3249_pp0_iter53_reg;
            p_read_61_reg_3249_pp0_iter55_reg <= p_read_61_reg_3249_pp0_iter54_reg;
            p_read_61_reg_3249_pp0_iter56_reg <= p_read_61_reg_3249_pp0_iter55_reg;
            p_read_61_reg_3249_pp0_iter57_reg <= p_read_61_reg_3249_pp0_iter56_reg;
            p_read_61_reg_3249_pp0_iter58_reg <= p_read_61_reg_3249_pp0_iter57_reg;
            p_read_61_reg_3249_pp0_iter59_reg <= p_read_61_reg_3249_pp0_iter58_reg;
            p_read_61_reg_3249_pp0_iter5_reg <= p_read_61_reg_3249_pp0_iter4_reg;
            p_read_61_reg_3249_pp0_iter60_reg <= p_read_61_reg_3249_pp0_iter59_reg;
            p_read_61_reg_3249_pp0_iter61_reg <= p_read_61_reg_3249_pp0_iter60_reg;
            p_read_61_reg_3249_pp0_iter62_reg <= p_read_61_reg_3249_pp0_iter61_reg;
            p_read_61_reg_3249_pp0_iter63_reg <= p_read_61_reg_3249_pp0_iter62_reg;
            p_read_61_reg_3249_pp0_iter64_reg <= p_read_61_reg_3249_pp0_iter63_reg;
            p_read_61_reg_3249_pp0_iter65_reg <= p_read_61_reg_3249_pp0_iter64_reg;
            p_read_61_reg_3249_pp0_iter66_reg <= p_read_61_reg_3249_pp0_iter65_reg;
            p_read_61_reg_3249_pp0_iter67_reg <= p_read_61_reg_3249_pp0_iter66_reg;
            p_read_61_reg_3249_pp0_iter68_reg <= p_read_61_reg_3249_pp0_iter67_reg;
            p_read_61_reg_3249_pp0_iter69_reg <= p_read_61_reg_3249_pp0_iter68_reg;
            p_read_61_reg_3249_pp0_iter6_reg <= p_read_61_reg_3249_pp0_iter5_reg;
            p_read_61_reg_3249_pp0_iter70_reg <= p_read_61_reg_3249_pp0_iter69_reg;
            p_read_61_reg_3249_pp0_iter71_reg <= p_read_61_reg_3249_pp0_iter70_reg;
            p_read_61_reg_3249_pp0_iter72_reg <= p_read_61_reg_3249_pp0_iter71_reg;
            p_read_61_reg_3249_pp0_iter73_reg <= p_read_61_reg_3249_pp0_iter72_reg;
            p_read_61_reg_3249_pp0_iter74_reg <= p_read_61_reg_3249_pp0_iter73_reg;
            p_read_61_reg_3249_pp0_iter75_reg <= p_read_61_reg_3249_pp0_iter74_reg;
            p_read_61_reg_3249_pp0_iter76_reg <= p_read_61_reg_3249_pp0_iter75_reg;
            p_read_61_reg_3249_pp0_iter7_reg <= p_read_61_reg_3249_pp0_iter6_reg;
            p_read_61_reg_3249_pp0_iter8_reg <= p_read_61_reg_3249_pp0_iter7_reg;
            p_read_61_reg_3249_pp0_iter9_reg <= p_read_61_reg_3249_pp0_iter8_reg;
            p_read_62_reg_3254 <= p_read2_int_reg;
            p_read_62_reg_3254_pp0_iter10_reg <= p_read_62_reg_3254_pp0_iter9_reg;
            p_read_62_reg_3254_pp0_iter11_reg <= p_read_62_reg_3254_pp0_iter10_reg;
            p_read_62_reg_3254_pp0_iter12_reg <= p_read_62_reg_3254_pp0_iter11_reg;
            p_read_62_reg_3254_pp0_iter13_reg <= p_read_62_reg_3254_pp0_iter12_reg;
            p_read_62_reg_3254_pp0_iter14_reg <= p_read_62_reg_3254_pp0_iter13_reg;
            p_read_62_reg_3254_pp0_iter15_reg <= p_read_62_reg_3254_pp0_iter14_reg;
            p_read_62_reg_3254_pp0_iter16_reg <= p_read_62_reg_3254_pp0_iter15_reg;
            p_read_62_reg_3254_pp0_iter17_reg <= p_read_62_reg_3254_pp0_iter16_reg;
            p_read_62_reg_3254_pp0_iter18_reg <= p_read_62_reg_3254_pp0_iter17_reg;
            p_read_62_reg_3254_pp0_iter19_reg <= p_read_62_reg_3254_pp0_iter18_reg;
            p_read_62_reg_3254_pp0_iter1_reg <= p_read_62_reg_3254;
            p_read_62_reg_3254_pp0_iter20_reg <= p_read_62_reg_3254_pp0_iter19_reg;
            p_read_62_reg_3254_pp0_iter21_reg <= p_read_62_reg_3254_pp0_iter20_reg;
            p_read_62_reg_3254_pp0_iter22_reg <= p_read_62_reg_3254_pp0_iter21_reg;
            p_read_62_reg_3254_pp0_iter23_reg <= p_read_62_reg_3254_pp0_iter22_reg;
            p_read_62_reg_3254_pp0_iter24_reg <= p_read_62_reg_3254_pp0_iter23_reg;
            p_read_62_reg_3254_pp0_iter25_reg <= p_read_62_reg_3254_pp0_iter24_reg;
            p_read_62_reg_3254_pp0_iter26_reg <= p_read_62_reg_3254_pp0_iter25_reg;
            p_read_62_reg_3254_pp0_iter27_reg <= p_read_62_reg_3254_pp0_iter26_reg;
            p_read_62_reg_3254_pp0_iter28_reg <= p_read_62_reg_3254_pp0_iter27_reg;
            p_read_62_reg_3254_pp0_iter29_reg <= p_read_62_reg_3254_pp0_iter28_reg;
            p_read_62_reg_3254_pp0_iter2_reg <= p_read_62_reg_3254_pp0_iter1_reg;
            p_read_62_reg_3254_pp0_iter30_reg <= p_read_62_reg_3254_pp0_iter29_reg;
            p_read_62_reg_3254_pp0_iter31_reg <= p_read_62_reg_3254_pp0_iter30_reg;
            p_read_62_reg_3254_pp0_iter32_reg <= p_read_62_reg_3254_pp0_iter31_reg;
            p_read_62_reg_3254_pp0_iter33_reg <= p_read_62_reg_3254_pp0_iter32_reg;
            p_read_62_reg_3254_pp0_iter34_reg <= p_read_62_reg_3254_pp0_iter33_reg;
            p_read_62_reg_3254_pp0_iter35_reg <= p_read_62_reg_3254_pp0_iter34_reg;
            p_read_62_reg_3254_pp0_iter36_reg <= p_read_62_reg_3254_pp0_iter35_reg;
            p_read_62_reg_3254_pp0_iter37_reg <= p_read_62_reg_3254_pp0_iter36_reg;
            p_read_62_reg_3254_pp0_iter38_reg <= p_read_62_reg_3254_pp0_iter37_reg;
            p_read_62_reg_3254_pp0_iter39_reg <= p_read_62_reg_3254_pp0_iter38_reg;
            p_read_62_reg_3254_pp0_iter3_reg <= p_read_62_reg_3254_pp0_iter2_reg;
            p_read_62_reg_3254_pp0_iter40_reg <= p_read_62_reg_3254_pp0_iter39_reg;
            p_read_62_reg_3254_pp0_iter41_reg <= p_read_62_reg_3254_pp0_iter40_reg;
            p_read_62_reg_3254_pp0_iter42_reg <= p_read_62_reg_3254_pp0_iter41_reg;
            p_read_62_reg_3254_pp0_iter43_reg <= p_read_62_reg_3254_pp0_iter42_reg;
            p_read_62_reg_3254_pp0_iter44_reg <= p_read_62_reg_3254_pp0_iter43_reg;
            p_read_62_reg_3254_pp0_iter45_reg <= p_read_62_reg_3254_pp0_iter44_reg;
            p_read_62_reg_3254_pp0_iter46_reg <= p_read_62_reg_3254_pp0_iter45_reg;
            p_read_62_reg_3254_pp0_iter47_reg <= p_read_62_reg_3254_pp0_iter46_reg;
            p_read_62_reg_3254_pp0_iter48_reg <= p_read_62_reg_3254_pp0_iter47_reg;
            p_read_62_reg_3254_pp0_iter49_reg <= p_read_62_reg_3254_pp0_iter48_reg;
            p_read_62_reg_3254_pp0_iter4_reg <= p_read_62_reg_3254_pp0_iter3_reg;
            p_read_62_reg_3254_pp0_iter50_reg <= p_read_62_reg_3254_pp0_iter49_reg;
            p_read_62_reg_3254_pp0_iter51_reg <= p_read_62_reg_3254_pp0_iter50_reg;
            p_read_62_reg_3254_pp0_iter52_reg <= p_read_62_reg_3254_pp0_iter51_reg;
            p_read_62_reg_3254_pp0_iter53_reg <= p_read_62_reg_3254_pp0_iter52_reg;
            p_read_62_reg_3254_pp0_iter54_reg <= p_read_62_reg_3254_pp0_iter53_reg;
            p_read_62_reg_3254_pp0_iter55_reg <= p_read_62_reg_3254_pp0_iter54_reg;
            p_read_62_reg_3254_pp0_iter56_reg <= p_read_62_reg_3254_pp0_iter55_reg;
            p_read_62_reg_3254_pp0_iter57_reg <= p_read_62_reg_3254_pp0_iter56_reg;
            p_read_62_reg_3254_pp0_iter58_reg <= p_read_62_reg_3254_pp0_iter57_reg;
            p_read_62_reg_3254_pp0_iter59_reg <= p_read_62_reg_3254_pp0_iter58_reg;
            p_read_62_reg_3254_pp0_iter5_reg <= p_read_62_reg_3254_pp0_iter4_reg;
            p_read_62_reg_3254_pp0_iter60_reg <= p_read_62_reg_3254_pp0_iter59_reg;
            p_read_62_reg_3254_pp0_iter61_reg <= p_read_62_reg_3254_pp0_iter60_reg;
            p_read_62_reg_3254_pp0_iter62_reg <= p_read_62_reg_3254_pp0_iter61_reg;
            p_read_62_reg_3254_pp0_iter63_reg <= p_read_62_reg_3254_pp0_iter62_reg;
            p_read_62_reg_3254_pp0_iter64_reg <= p_read_62_reg_3254_pp0_iter63_reg;
            p_read_62_reg_3254_pp0_iter65_reg <= p_read_62_reg_3254_pp0_iter64_reg;
            p_read_62_reg_3254_pp0_iter66_reg <= p_read_62_reg_3254_pp0_iter65_reg;
            p_read_62_reg_3254_pp0_iter67_reg <= p_read_62_reg_3254_pp0_iter66_reg;
            p_read_62_reg_3254_pp0_iter68_reg <= p_read_62_reg_3254_pp0_iter67_reg;
            p_read_62_reg_3254_pp0_iter69_reg <= p_read_62_reg_3254_pp0_iter68_reg;
            p_read_62_reg_3254_pp0_iter6_reg <= p_read_62_reg_3254_pp0_iter5_reg;
            p_read_62_reg_3254_pp0_iter70_reg <= p_read_62_reg_3254_pp0_iter69_reg;
            p_read_62_reg_3254_pp0_iter71_reg <= p_read_62_reg_3254_pp0_iter70_reg;
            p_read_62_reg_3254_pp0_iter72_reg <= p_read_62_reg_3254_pp0_iter71_reg;
            p_read_62_reg_3254_pp0_iter73_reg <= p_read_62_reg_3254_pp0_iter72_reg;
            p_read_62_reg_3254_pp0_iter74_reg <= p_read_62_reg_3254_pp0_iter73_reg;
            p_read_62_reg_3254_pp0_iter75_reg <= p_read_62_reg_3254_pp0_iter74_reg;
            p_read_62_reg_3254_pp0_iter76_reg <= p_read_62_reg_3254_pp0_iter75_reg;
            p_read_62_reg_3254_pp0_iter7_reg <= p_read_62_reg_3254_pp0_iter6_reg;
            p_read_62_reg_3254_pp0_iter8_reg <= p_read_62_reg_3254_pp0_iter7_reg;
            p_read_62_reg_3254_pp0_iter9_reg <= p_read_62_reg_3254_pp0_iter8_reg;
            p_read_63_reg_3259 <= p_read1_int_reg;
            p_read_63_reg_3259_pp0_iter10_reg <= p_read_63_reg_3259_pp0_iter9_reg;
            p_read_63_reg_3259_pp0_iter11_reg <= p_read_63_reg_3259_pp0_iter10_reg;
            p_read_63_reg_3259_pp0_iter12_reg <= p_read_63_reg_3259_pp0_iter11_reg;
            p_read_63_reg_3259_pp0_iter13_reg <= p_read_63_reg_3259_pp0_iter12_reg;
            p_read_63_reg_3259_pp0_iter14_reg <= p_read_63_reg_3259_pp0_iter13_reg;
            p_read_63_reg_3259_pp0_iter15_reg <= p_read_63_reg_3259_pp0_iter14_reg;
            p_read_63_reg_3259_pp0_iter16_reg <= p_read_63_reg_3259_pp0_iter15_reg;
            p_read_63_reg_3259_pp0_iter17_reg <= p_read_63_reg_3259_pp0_iter16_reg;
            p_read_63_reg_3259_pp0_iter18_reg <= p_read_63_reg_3259_pp0_iter17_reg;
            p_read_63_reg_3259_pp0_iter19_reg <= p_read_63_reg_3259_pp0_iter18_reg;
            p_read_63_reg_3259_pp0_iter1_reg <= p_read_63_reg_3259;
            p_read_63_reg_3259_pp0_iter20_reg <= p_read_63_reg_3259_pp0_iter19_reg;
            p_read_63_reg_3259_pp0_iter21_reg <= p_read_63_reg_3259_pp0_iter20_reg;
            p_read_63_reg_3259_pp0_iter22_reg <= p_read_63_reg_3259_pp0_iter21_reg;
            p_read_63_reg_3259_pp0_iter23_reg <= p_read_63_reg_3259_pp0_iter22_reg;
            p_read_63_reg_3259_pp0_iter24_reg <= p_read_63_reg_3259_pp0_iter23_reg;
            p_read_63_reg_3259_pp0_iter25_reg <= p_read_63_reg_3259_pp0_iter24_reg;
            p_read_63_reg_3259_pp0_iter26_reg <= p_read_63_reg_3259_pp0_iter25_reg;
            p_read_63_reg_3259_pp0_iter27_reg <= p_read_63_reg_3259_pp0_iter26_reg;
            p_read_63_reg_3259_pp0_iter28_reg <= p_read_63_reg_3259_pp0_iter27_reg;
            p_read_63_reg_3259_pp0_iter29_reg <= p_read_63_reg_3259_pp0_iter28_reg;
            p_read_63_reg_3259_pp0_iter2_reg <= p_read_63_reg_3259_pp0_iter1_reg;
            p_read_63_reg_3259_pp0_iter30_reg <= p_read_63_reg_3259_pp0_iter29_reg;
            p_read_63_reg_3259_pp0_iter31_reg <= p_read_63_reg_3259_pp0_iter30_reg;
            p_read_63_reg_3259_pp0_iter32_reg <= p_read_63_reg_3259_pp0_iter31_reg;
            p_read_63_reg_3259_pp0_iter33_reg <= p_read_63_reg_3259_pp0_iter32_reg;
            p_read_63_reg_3259_pp0_iter34_reg <= p_read_63_reg_3259_pp0_iter33_reg;
            p_read_63_reg_3259_pp0_iter35_reg <= p_read_63_reg_3259_pp0_iter34_reg;
            p_read_63_reg_3259_pp0_iter36_reg <= p_read_63_reg_3259_pp0_iter35_reg;
            p_read_63_reg_3259_pp0_iter37_reg <= p_read_63_reg_3259_pp0_iter36_reg;
            p_read_63_reg_3259_pp0_iter38_reg <= p_read_63_reg_3259_pp0_iter37_reg;
            p_read_63_reg_3259_pp0_iter39_reg <= p_read_63_reg_3259_pp0_iter38_reg;
            p_read_63_reg_3259_pp0_iter3_reg <= p_read_63_reg_3259_pp0_iter2_reg;
            p_read_63_reg_3259_pp0_iter40_reg <= p_read_63_reg_3259_pp0_iter39_reg;
            p_read_63_reg_3259_pp0_iter41_reg <= p_read_63_reg_3259_pp0_iter40_reg;
            p_read_63_reg_3259_pp0_iter42_reg <= p_read_63_reg_3259_pp0_iter41_reg;
            p_read_63_reg_3259_pp0_iter43_reg <= p_read_63_reg_3259_pp0_iter42_reg;
            p_read_63_reg_3259_pp0_iter44_reg <= p_read_63_reg_3259_pp0_iter43_reg;
            p_read_63_reg_3259_pp0_iter45_reg <= p_read_63_reg_3259_pp0_iter44_reg;
            p_read_63_reg_3259_pp0_iter46_reg <= p_read_63_reg_3259_pp0_iter45_reg;
            p_read_63_reg_3259_pp0_iter47_reg <= p_read_63_reg_3259_pp0_iter46_reg;
            p_read_63_reg_3259_pp0_iter48_reg <= p_read_63_reg_3259_pp0_iter47_reg;
            p_read_63_reg_3259_pp0_iter49_reg <= p_read_63_reg_3259_pp0_iter48_reg;
            p_read_63_reg_3259_pp0_iter4_reg <= p_read_63_reg_3259_pp0_iter3_reg;
            p_read_63_reg_3259_pp0_iter50_reg <= p_read_63_reg_3259_pp0_iter49_reg;
            p_read_63_reg_3259_pp0_iter51_reg <= p_read_63_reg_3259_pp0_iter50_reg;
            p_read_63_reg_3259_pp0_iter52_reg <= p_read_63_reg_3259_pp0_iter51_reg;
            p_read_63_reg_3259_pp0_iter53_reg <= p_read_63_reg_3259_pp0_iter52_reg;
            p_read_63_reg_3259_pp0_iter54_reg <= p_read_63_reg_3259_pp0_iter53_reg;
            p_read_63_reg_3259_pp0_iter55_reg <= p_read_63_reg_3259_pp0_iter54_reg;
            p_read_63_reg_3259_pp0_iter56_reg <= p_read_63_reg_3259_pp0_iter55_reg;
            p_read_63_reg_3259_pp0_iter57_reg <= p_read_63_reg_3259_pp0_iter56_reg;
            p_read_63_reg_3259_pp0_iter58_reg <= p_read_63_reg_3259_pp0_iter57_reg;
            p_read_63_reg_3259_pp0_iter59_reg <= p_read_63_reg_3259_pp0_iter58_reg;
            p_read_63_reg_3259_pp0_iter5_reg <= p_read_63_reg_3259_pp0_iter4_reg;
            p_read_63_reg_3259_pp0_iter60_reg <= p_read_63_reg_3259_pp0_iter59_reg;
            p_read_63_reg_3259_pp0_iter61_reg <= p_read_63_reg_3259_pp0_iter60_reg;
            p_read_63_reg_3259_pp0_iter62_reg <= p_read_63_reg_3259_pp0_iter61_reg;
            p_read_63_reg_3259_pp0_iter63_reg <= p_read_63_reg_3259_pp0_iter62_reg;
            p_read_63_reg_3259_pp0_iter64_reg <= p_read_63_reg_3259_pp0_iter63_reg;
            p_read_63_reg_3259_pp0_iter65_reg <= p_read_63_reg_3259_pp0_iter64_reg;
            p_read_63_reg_3259_pp0_iter66_reg <= p_read_63_reg_3259_pp0_iter65_reg;
            p_read_63_reg_3259_pp0_iter67_reg <= p_read_63_reg_3259_pp0_iter66_reg;
            p_read_63_reg_3259_pp0_iter68_reg <= p_read_63_reg_3259_pp0_iter67_reg;
            p_read_63_reg_3259_pp0_iter69_reg <= p_read_63_reg_3259_pp0_iter68_reg;
            p_read_63_reg_3259_pp0_iter6_reg <= p_read_63_reg_3259_pp0_iter5_reg;
            p_read_63_reg_3259_pp0_iter70_reg <= p_read_63_reg_3259_pp0_iter69_reg;
            p_read_63_reg_3259_pp0_iter71_reg <= p_read_63_reg_3259_pp0_iter70_reg;
            p_read_63_reg_3259_pp0_iter72_reg <= p_read_63_reg_3259_pp0_iter71_reg;
            p_read_63_reg_3259_pp0_iter73_reg <= p_read_63_reg_3259_pp0_iter72_reg;
            p_read_63_reg_3259_pp0_iter74_reg <= p_read_63_reg_3259_pp0_iter73_reg;
            p_read_63_reg_3259_pp0_iter75_reg <= p_read_63_reg_3259_pp0_iter74_reg;
            p_read_63_reg_3259_pp0_iter76_reg <= p_read_63_reg_3259_pp0_iter75_reg;
            p_read_63_reg_3259_pp0_iter7_reg <= p_read_63_reg_3259_pp0_iter6_reg;
            p_read_63_reg_3259_pp0_iter8_reg <= p_read_63_reg_3259_pp0_iter7_reg;
            p_read_63_reg_3259_pp0_iter9_reg <= p_read_63_reg_3259_pp0_iter8_reg;
            x_read_reg_3281 <= x_int_reg;
            x_read_reg_3281_pp0_iter10_reg <= x_read_reg_3281_pp0_iter9_reg;
            x_read_reg_3281_pp0_iter11_reg <= x_read_reg_3281_pp0_iter10_reg;
            x_read_reg_3281_pp0_iter12_reg <= x_read_reg_3281_pp0_iter11_reg;
            x_read_reg_3281_pp0_iter13_reg <= x_read_reg_3281_pp0_iter12_reg;
            x_read_reg_3281_pp0_iter14_reg <= x_read_reg_3281_pp0_iter13_reg;
            x_read_reg_3281_pp0_iter15_reg <= x_read_reg_3281_pp0_iter14_reg;
            x_read_reg_3281_pp0_iter16_reg <= x_read_reg_3281_pp0_iter15_reg;
            x_read_reg_3281_pp0_iter17_reg <= x_read_reg_3281_pp0_iter16_reg;
            x_read_reg_3281_pp0_iter18_reg <= x_read_reg_3281_pp0_iter17_reg;
            x_read_reg_3281_pp0_iter19_reg <= x_read_reg_3281_pp0_iter18_reg;
            x_read_reg_3281_pp0_iter1_reg <= x_read_reg_3281;
            x_read_reg_3281_pp0_iter20_reg <= x_read_reg_3281_pp0_iter19_reg;
            x_read_reg_3281_pp0_iter2_reg <= x_read_reg_3281_pp0_iter1_reg;
            x_read_reg_3281_pp0_iter3_reg <= x_read_reg_3281_pp0_iter2_reg;
            x_read_reg_3281_pp0_iter4_reg <= x_read_reg_3281_pp0_iter3_reg;
            x_read_reg_3281_pp0_iter5_reg <= x_read_reg_3281_pp0_iter4_reg;
            x_read_reg_3281_pp0_iter6_reg <= x_read_reg_3281_pp0_iter5_reg;
            x_read_reg_3281_pp0_iter7_reg <= x_read_reg_3281_pp0_iter6_reg;
            x_read_reg_3281_pp0_iter8_reg <= x_read_reg_3281_pp0_iter7_reg;
            x_read_reg_3281_pp0_iter9_reg <= x_read_reg_3281_pp0_iter8_reg;
            y_read_reg_3275 <= y_int_reg;
            y_read_reg_3275_pp0_iter10_reg <= y_read_reg_3275_pp0_iter9_reg;
            y_read_reg_3275_pp0_iter11_reg <= y_read_reg_3275_pp0_iter10_reg;
            y_read_reg_3275_pp0_iter12_reg <= y_read_reg_3275_pp0_iter11_reg;
            y_read_reg_3275_pp0_iter13_reg <= y_read_reg_3275_pp0_iter12_reg;
            y_read_reg_3275_pp0_iter14_reg <= y_read_reg_3275_pp0_iter13_reg;
            y_read_reg_3275_pp0_iter15_reg <= y_read_reg_3275_pp0_iter14_reg;
            y_read_reg_3275_pp0_iter16_reg <= y_read_reg_3275_pp0_iter15_reg;
            y_read_reg_3275_pp0_iter17_reg <= y_read_reg_3275_pp0_iter16_reg;
            y_read_reg_3275_pp0_iter18_reg <= y_read_reg_3275_pp0_iter17_reg;
            y_read_reg_3275_pp0_iter19_reg <= y_read_reg_3275_pp0_iter18_reg;
            y_read_reg_3275_pp0_iter1_reg <= y_read_reg_3275;
            y_read_reg_3275_pp0_iter20_reg <= y_read_reg_3275_pp0_iter19_reg;
            y_read_reg_3275_pp0_iter2_reg <= y_read_reg_3275_pp0_iter1_reg;
            y_read_reg_3275_pp0_iter3_reg <= y_read_reg_3275_pp0_iter2_reg;
            y_read_reg_3275_pp0_iter4_reg <= y_read_reg_3275_pp0_iter3_reg;
            y_read_reg_3275_pp0_iter5_reg <= y_read_reg_3275_pp0_iter4_reg;
            y_read_reg_3275_pp0_iter6_reg <= y_read_reg_3275_pp0_iter5_reg;
            y_read_reg_3275_pp0_iter7_reg <= y_read_reg_3275_pp0_iter6_reg;
            y_read_reg_3275_pp0_iter8_reg <= y_read_reg_3275_pp0_iter7_reg;
            y_read_reg_3275_pp0_iter9_reg <= y_read_reg_3275_pp0_iter8_reg;
            z_read_reg_3269 <= z_int_reg;
            z_read_reg_3269_pp0_iter10_reg <= z_read_reg_3269_pp0_iter9_reg;
            z_read_reg_3269_pp0_iter11_reg <= z_read_reg_3269_pp0_iter10_reg;
            z_read_reg_3269_pp0_iter12_reg <= z_read_reg_3269_pp0_iter11_reg;
            z_read_reg_3269_pp0_iter13_reg <= z_read_reg_3269_pp0_iter12_reg;
            z_read_reg_3269_pp0_iter14_reg <= z_read_reg_3269_pp0_iter13_reg;
            z_read_reg_3269_pp0_iter15_reg <= z_read_reg_3269_pp0_iter14_reg;
            z_read_reg_3269_pp0_iter16_reg <= z_read_reg_3269_pp0_iter15_reg;
            z_read_reg_3269_pp0_iter17_reg <= z_read_reg_3269_pp0_iter16_reg;
            z_read_reg_3269_pp0_iter18_reg <= z_read_reg_3269_pp0_iter17_reg;
            z_read_reg_3269_pp0_iter19_reg <= z_read_reg_3269_pp0_iter18_reg;
            z_read_reg_3269_pp0_iter1_reg <= z_read_reg_3269;
            z_read_reg_3269_pp0_iter20_reg <= z_read_reg_3269_pp0_iter19_reg;
            z_read_reg_3269_pp0_iter2_reg <= z_read_reg_3269_pp0_iter1_reg;
            z_read_reg_3269_pp0_iter3_reg <= z_read_reg_3269_pp0_iter2_reg;
            z_read_reg_3269_pp0_iter4_reg <= z_read_reg_3269_pp0_iter3_reg;
            z_read_reg_3269_pp0_iter5_reg <= z_read_reg_3269_pp0_iter4_reg;
            z_read_reg_3269_pp0_iter6_reg <= z_read_reg_3269_pp0_iter5_reg;
            z_read_reg_3269_pp0_iter7_reg <= z_read_reg_3269_pp0_iter6_reg;
            z_read_reg_3269_pp0_iter8_reg <= z_read_reg_3269_pp0_iter7_reg;
            z_read_reg_3269_pp0_iter9_reg <= z_read_reg_3269_pp0_iter8_reg;
        end
    end

    assign H_offset_read_read_fu_158_p2 = H_offset_int_reg;

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_phi_reg_pp0_iter0_phi_ln112_10_reg_1568 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_11_reg_1583 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_12_reg_1598 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_13_reg_1613 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_14_reg_1628 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_15_reg_1643 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_1_reg_1673 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_2_reg_1688 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_3_reg_1703 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_4_reg_1478 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_5_reg_1493 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_6_reg_1508 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_7_reg_1523 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_8_reg_1538 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_9_reg_1553 = 'bx;

    assign ap_phi_reg_pp0_iter0_phi_ln112_reg_1658 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag101_0_reg_1212 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag104_0_reg_1193 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag107_0_reg_1174 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag110_0_reg_1307 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag113_0_reg_1288 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag116_0_reg_1269 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag119_0_reg_1250 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag11_0_reg_566 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag122_0_reg_1383 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag125_0_reg_1345 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag128_0_reg_1326 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag131_0_reg_1364 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag134_0_reg_1402 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag137_0_reg_1421 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag140_0_reg_1440 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag143_0_reg_1459 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag14_0_reg_699 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag17_0_reg_680 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag20_0_reg_661 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag23_0_reg_642 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag26_0_reg_775 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag29_0_reg_756 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag32_0_reg_718 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag35_0_reg_737 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag38_0_reg_794 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag41_0_reg_813 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag44_0_reg_832 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag47_0_reg_851 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag4_0_reg_604 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag50_0_reg_870 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag53_0_reg_889 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag56_0_reg_908 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag59_0_reg_927 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag62_0_reg_946 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag65_0_reg_965 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag68_0_reg_984 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag71_0_reg_1003 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag74_0_reg_1022 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag77_0_reg_1041 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag80_0_reg_1060 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag83_0_reg_1079 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag86_0_reg_1098 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag89_0_reg_1117 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag8_0_reg_585 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag92_0_reg_1136 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag95_0_reg_1155 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag98_0_reg_1231 = 'bx;

    assign ap_phi_reg_pp0_iter0_write_flag_0_reg_623 = 'bx;

    assign ap_return_0 = select_ln112_fu_2242_p3;

    assign ap_return_1 = select_ln112_1_fu_2248_p3;

    assign ap_return_10 = select_ln112_10_fu_2302_p3;

    assign ap_return_11 = select_ln112_11_fu_2308_p3;

    assign ap_return_12 = select_ln112_12_fu_2314_p3;

    assign ap_return_13 = select_ln112_13_fu_2320_p3;

    assign ap_return_14 = select_ln112_14_fu_2326_p3;

    assign ap_return_15 = select_ln112_15_fu_2332_p3;

    assign ap_return_16 = select_ln112_16_fu_2338_p3;

    assign ap_return_17 = select_ln112_17_fu_2344_p3;

    assign ap_return_18 = select_ln112_18_fu_2350_p3;

    assign ap_return_19 = select_ln112_19_fu_2356_p3;

    assign ap_return_2 = select_ln112_2_fu_2254_p3;

    assign ap_return_20 = select_ln112_20_fu_2362_p3;

    assign ap_return_21 = select_ln112_21_fu_2368_p3;

    assign ap_return_22 = select_ln112_22_fu_2374_p3;

    assign ap_return_23 = select_ln112_23_fu_2380_p3;

    assign ap_return_24 = select_ln112_24_fu_2386_p3;

    assign ap_return_25 = select_ln112_25_fu_2392_p3;

    assign ap_return_26 = select_ln112_26_fu_2398_p3;

    assign ap_return_27 = select_ln112_27_fu_2404_p3;

    assign ap_return_28 = select_ln112_28_fu_2410_p3;

    assign ap_return_29 = select_ln112_29_fu_2416_p3;

    assign ap_return_3 = select_ln112_3_fu_2260_p3;

    assign ap_return_30 = select_ln112_30_fu_2422_p3;

    assign ap_return_31 = select_ln112_31_fu_2428_p3;

    assign ap_return_32 = select_ln112_32_fu_2434_p3;

    assign ap_return_33 = select_ln112_33_fu_2440_p3;

    assign ap_return_34 = select_ln112_34_fu_2446_p3;

    assign ap_return_35 = select_ln112_35_fu_2452_p3;

    assign ap_return_36 = select_ln112_36_fu_2458_p3;

    assign ap_return_37 = select_ln112_37_fu_2464_p3;

    assign ap_return_38 = select_ln112_38_fu_2470_p3;

    assign ap_return_39 = select_ln112_39_fu_2476_p3;

    assign ap_return_4 = select_ln112_4_fu_2266_p3;

    assign ap_return_40 = select_ln112_40_fu_2482_p3;

    assign ap_return_41 = select_ln112_41_fu_2488_p3;

    assign ap_return_42 = select_ln112_42_fu_2494_p3;

    assign ap_return_43 = select_ln112_43_fu_2500_p3;

    assign ap_return_44 = select_ln112_44_fu_2506_p3;

    assign ap_return_45 = select_ln112_45_fu_2512_p3;

    assign ap_return_46 = select_ln112_46_fu_2518_p3;

    assign ap_return_47 = select_ln112_47_fu_2524_p3;

    assign ap_return_48 = ap_phi_reg_pp0_iter77_phi_ln112_4_reg_1478;

    assign ap_return_49 = ap_phi_reg_pp0_iter77_phi_ln112_5_reg_1493;

    assign ap_return_5 = select_ln112_5_fu_2272_p3;

    assign ap_return_50 = ap_phi_reg_pp0_iter77_phi_ln112_6_reg_1508;

    assign ap_return_51 = ap_phi_reg_pp0_iter77_phi_ln112_7_reg_1523;

    assign ap_return_52 = ap_phi_reg_pp0_iter77_phi_ln112_8_reg_1538;

    assign ap_return_53 = ap_phi_reg_pp0_iter77_phi_ln112_9_reg_1553;

    assign ap_return_54 = ap_phi_reg_pp0_iter77_phi_ln112_10_reg_1568;

    assign ap_return_55 = ap_phi_reg_pp0_iter77_phi_ln112_11_reg_1583;

    assign ap_return_56 = ap_phi_reg_pp0_iter77_phi_ln112_12_reg_1598;

    assign ap_return_57 = ap_phi_reg_pp0_iter77_phi_ln112_13_reg_1613;

    assign ap_return_58 = ap_phi_reg_pp0_iter77_phi_ln112_14_reg_1628;

    assign ap_return_59 = ap_phi_reg_pp0_iter77_phi_ln112_15_reg_1643;

    assign ap_return_6 = select_ln112_6_fu_2278_p3;

    assign ap_return_60 = ap_phi_reg_pp0_iter77_phi_ln112_reg_1658;

    assign ap_return_61 = ap_phi_reg_pp0_iter77_phi_ln112_1_reg_1673;

    assign ap_return_62 = ap_phi_reg_pp0_iter77_phi_ln112_2_reg_1688;

    assign ap_return_63 = ap_phi_reg_pp0_iter77_phi_ln112_3_reg_1703;

    assign ap_return_7 = select_ln112_7_fu_2284_p3;

    assign ap_return_8 = select_ln112_8_fu_2290_p3;

    assign ap_return_9 = select_ln112_9_fu_2296_p3;

    assign select_ln112_10_fu_2302_p3 = ((ap_phi_reg_pp0_iter77_write_flag32_0_reg_718[0:0] == 1'b1) ? H_0_27_reg_3908 : p_read_54_reg_3214_pp0_iter76_reg);

    assign select_ln112_11_fu_2308_p3 = ((ap_phi_reg_pp0_iter77_write_flag35_0_reg_737[0:0] == 1'b1) ? H_0_27_reg_3908 : p_read_53_reg_3209_pp0_iter76_reg);

    assign select_ln112_12_fu_2314_p3 = ((ap_phi_reg_pp0_iter77_write_flag38_0_reg_794[0:0] == 1'b1) ? H_0_3_reg_3916 : p_read_52_reg_3204_pp0_iter76_reg);

    assign select_ln112_13_fu_2320_p3 = ((ap_phi_reg_pp0_iter77_write_flag41_0_reg_813[0:0] == 1'b1) ? H_0_3_reg_3916 : p_read_51_reg_3199_pp0_iter76_reg);

    assign select_ln112_14_fu_2326_p3 = ((ap_phi_reg_pp0_iter77_write_flag44_0_reg_832[0:0] == 1'b1) ? H_0_3_reg_3916 : p_read_50_reg_3194_pp0_iter76_reg);

    assign select_ln112_15_fu_2332_p3 = ((ap_phi_reg_pp0_iter77_write_flag47_0_reg_851[0:0] == 1'b1) ? H_0_3_reg_3916 : p_read_49_reg_3189_pp0_iter76_reg);

    assign select_ln112_16_fu_2338_p3 = ((ap_phi_reg_pp0_iter77_write_flag50_0_reg_870[0:0] == 1'b1) ? H_1_0_reg_3924 : p_read_48_reg_3184_pp0_iter76_reg);

    assign select_ln112_17_fu_2344_p3 = ((ap_phi_reg_pp0_iter77_write_flag53_0_reg_889[0:0] == 1'b1) ? H_1_0_reg_3924 : p_read_47_reg_3179_pp0_iter76_reg);

    assign select_ln112_18_fu_2350_p3 = ((ap_phi_reg_pp0_iter77_write_flag56_0_reg_908[0:0] == 1'b1) ? H_1_0_reg_3924 : p_read_46_reg_3174_pp0_iter76_reg);

    assign select_ln112_19_fu_2356_p3 = ((ap_phi_reg_pp0_iter77_write_flag59_0_reg_927[0:0] == 1'b1) ? H_1_0_reg_3924 : p_read_45_reg_3169_pp0_iter76_reg);

    assign select_ln112_1_fu_2248_p3 = ((ap_phi_reg_pp0_iter77_write_flag4_0_reg_604[0:0] == 1'b1) ? H_0_03_reg_3892 : p_read_63_reg_3259_pp0_iter76_reg);

    assign select_ln112_20_fu_2362_p3 = ((ap_phi_reg_pp0_iter77_write_flag62_0_reg_946[0:0] == 1'b1) ? H_1_1_reg_3932 : p_read_44_reg_3164_pp0_iter76_reg);

    assign select_ln112_21_fu_2368_p3 = ((ap_phi_reg_pp0_iter77_write_flag65_0_reg_965[0:0] == 1'b1) ? H_1_1_reg_3932 : p_read_43_reg_3159_pp0_iter76_reg);

    assign select_ln112_22_fu_2374_p3 = ((ap_phi_reg_pp0_iter77_write_flag68_0_reg_984[0:0] == 1'b1) ? H_1_1_reg_3932 : p_read_42_reg_3154_pp0_iter76_reg);

    assign select_ln112_23_fu_2380_p3 = ((ap_phi_reg_pp0_iter77_write_flag71_0_reg_1003[0:0] == 1'b1) ? H_1_1_reg_3932 : p_read_41_reg_3149_pp0_iter76_reg);

    assign select_ln112_24_fu_2386_p3 = ((ap_phi_reg_pp0_iter77_write_flag74_0_reg_1022[0:0] == 1'b1) ? H_1_2_reg_3940 : p_read_40_reg_3144_pp0_iter76_reg);

    assign select_ln112_25_fu_2392_p3 = ((ap_phi_reg_pp0_iter77_write_flag77_0_reg_1041[0:0] == 1'b1) ? H_1_2_reg_3940 : p_read_39_reg_3139_pp0_iter76_reg);

    assign select_ln112_26_fu_2398_p3 = ((ap_phi_reg_pp0_iter77_write_flag80_0_reg_1060[0:0] == 1'b1) ? H_1_2_reg_3940 : p_read_38_reg_3134_pp0_iter76_reg);

    assign select_ln112_27_fu_2404_p3 = ((ap_phi_reg_pp0_iter77_write_flag83_0_reg_1079[0:0] == 1'b1) ? H_1_2_reg_3940 : p_read_37_reg_3129_pp0_iter76_reg);

    assign select_ln112_28_fu_2410_p3 = ((ap_phi_reg_pp0_iter77_write_flag86_0_reg_1098[0:0] == 1'b1) ? H_1_3_reg_3948 : p_read_36_reg_3124_pp0_iter76_reg);

    assign select_ln112_29_fu_2416_p3 = ((ap_phi_reg_pp0_iter77_write_flag89_0_reg_1117[0:0] == 1'b1) ? H_1_3_reg_3948 : p_read_35_reg_3119_pp0_iter76_reg);

    assign select_ln112_2_fu_2254_p3 = ((ap_phi_reg_pp0_iter77_write_flag8_0_reg_585[0:0] == 1'b1) ? H_0_03_reg_3892 : p_read_62_reg_3254_pp0_iter76_reg);

    assign select_ln112_30_fu_2422_p3 = ((ap_phi_reg_pp0_iter77_write_flag92_0_reg_1136[0:0] == 1'b1) ? H_1_3_reg_3948 : p_read_34_reg_3114_pp0_iter76_reg);

    assign select_ln112_31_fu_2428_p3 = ((ap_phi_reg_pp0_iter77_write_flag95_0_reg_1155[0:0] == 1'b1) ? H_1_3_reg_3948 : p_read_33_reg_3109_pp0_iter76_reg);

    assign select_ln112_32_fu_2434_p3 = ((ap_phi_reg_pp0_iter77_write_flag98_0_reg_1231[0:0] == 1'b1) ? H_2_0_reg_3956 : p_read_32_reg_3104_pp0_iter76_reg);

    assign select_ln112_33_fu_2440_p3 = ((ap_phi_reg_pp0_iter77_write_flag101_0_reg_1212[0:0] == 1'b1) ? H_2_0_reg_3956 : p_read_31_reg_3099_pp0_iter76_reg);

    assign select_ln112_34_fu_2446_p3 = ((ap_phi_reg_pp0_iter77_write_flag104_0_reg_1193[0:0] == 1'b1) ? H_2_0_reg_3956 : p_read_30_reg_3094_pp0_iter76_reg);

    assign select_ln112_35_fu_2452_p3 = ((ap_phi_reg_pp0_iter77_write_flag107_0_reg_1174[0:0] == 1'b1) ? H_2_0_reg_3956 : p_read_29_reg_3089_pp0_iter76_reg);

    assign select_ln112_36_fu_2458_p3 = ((ap_phi_reg_pp0_iter77_write_flag110_0_reg_1307[0:0] == 1'b1) ? H_2_1_reg_3964 : p_read_28_reg_3084_pp0_iter76_reg);

    assign select_ln112_37_fu_2464_p3 = ((ap_phi_reg_pp0_iter77_write_flag113_0_reg_1288[0:0] == 1'b1) ? H_2_1_reg_3964 : p_read_27_reg_3079_pp0_iter76_reg);

    assign select_ln112_38_fu_2470_p3 = ((ap_phi_reg_pp0_iter77_write_flag116_0_reg_1269[0:0] == 1'b1) ? H_2_1_reg_3964 : p_read_26_reg_3074_pp0_iter76_reg);

    assign select_ln112_39_fu_2476_p3 = ((ap_phi_reg_pp0_iter77_write_flag119_0_reg_1250[0:0] == 1'b1) ? H_2_1_reg_3964 : p_read_25_reg_3069_pp0_iter76_reg);

    assign select_ln112_3_fu_2260_p3 = ((ap_phi_reg_pp0_iter77_write_flag11_0_reg_566[0:0] == 1'b1) ? H_0_03_reg_3892 : p_read_61_reg_3249_pp0_iter76_reg);

    assign select_ln112_40_fu_2482_p3 = ((ap_phi_reg_pp0_iter77_write_flag122_0_reg_1383[0:0] == 1'b1) ? H_2_2_reg_3972 : p_read_24_reg_3064_pp0_iter76_reg);

    assign select_ln112_41_fu_2488_p3 = ((ap_phi_reg_pp0_iter77_write_flag125_0_reg_1345[0:0] == 1'b1) ? H_2_2_reg_3972 : p_read_23_reg_3059_pp0_iter76_reg);

    assign select_ln112_42_fu_2494_p3 = ((ap_phi_reg_pp0_iter77_write_flag128_0_reg_1326[0:0] == 1'b1) ? H_2_2_reg_3972 : p_read_22_reg_3054_pp0_iter76_reg);

    assign select_ln112_43_fu_2500_p3 = ((ap_phi_reg_pp0_iter77_write_flag131_0_reg_1364[0:0] == 1'b1) ? H_2_2_reg_3972 : p_read_21_reg_3049_pp0_iter76_reg);

    assign select_ln112_44_fu_2506_p3 = ((ap_phi_reg_pp0_iter77_write_flag134_0_reg_1402[0:0] == 1'b1) ? H_2_3_reg_3980 : p_read_20_reg_3044_pp0_iter76_reg);

    assign select_ln112_45_fu_2512_p3 = ((ap_phi_reg_pp0_iter77_write_flag137_0_reg_1421[0:0] == 1'b1) ? H_2_3_reg_3980 : p_read_19_reg_3039_pp0_iter76_reg);

    assign select_ln112_46_fu_2518_p3 = ((ap_phi_reg_pp0_iter77_write_flag140_0_reg_1440[0:0] == 1'b1) ? H_2_3_reg_3980 : p_read_18_reg_3034_pp0_iter76_reg);

    assign select_ln112_47_fu_2524_p3 = ((ap_phi_reg_pp0_iter77_write_flag143_0_reg_1459[0:0] == 1'b1) ? H_2_3_reg_3980 : p_read_17_reg_3029_pp0_iter76_reg);

    assign select_ln112_4_fu_2266_p3 = ((ap_phi_reg_pp0_iter77_write_flag14_0_reg_699[0:0] == 1'b1) ? H_0_16_reg_3900 : p_read_60_reg_3244_pp0_iter76_reg);

    assign select_ln112_5_fu_2272_p3 = ((ap_phi_reg_pp0_iter77_write_flag17_0_reg_680[0:0] == 1'b1) ? H_0_16_reg_3900 : p_read_59_reg_3239_pp0_iter76_reg);

    assign select_ln112_6_fu_2278_p3 = ((ap_phi_reg_pp0_iter77_write_flag20_0_reg_661[0:0] == 1'b1) ? H_0_16_reg_3900 : p_read_58_reg_3234_pp0_iter76_reg);

    assign select_ln112_7_fu_2284_p3 = ((ap_phi_reg_pp0_iter77_write_flag23_0_reg_642[0:0] == 1'b1) ? H_0_16_reg_3900 : p_read_57_reg_3229_pp0_iter76_reg);

    assign select_ln112_8_fu_2290_p3 = ((ap_phi_reg_pp0_iter77_write_flag26_0_reg_775[0:0] == 1'b1) ? H_0_27_reg_3908 : p_read_56_reg_3224_pp0_iter76_reg);

    assign select_ln112_9_fu_2296_p3 = ((ap_phi_reg_pp0_iter77_write_flag29_0_reg_756[0:0] == 1'b1) ? H_0_27_reg_3908 : p_read_55_reg_3219_pp0_iter76_reg);

    assign select_ln112_fu_2242_p3 = ((ap_phi_reg_pp0_iter77_write_flag_0_reg_623[0:0] == 1'b1) ? H_0_03_reg_3892 : p_read64_reg_3264_pp0_iter76_reg);

endmodule  //main_rpyxyzToH_double_s
