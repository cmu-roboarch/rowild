/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_scaled_fixed2ieee_63_1_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    in_val,
    prescale,
    ap_return
);

    parameter ap_ST_fsm_state1 = 9'd1;
    parameter ap_ST_fsm_state2 = 9'd2;
    parameter ap_ST_fsm_state3 = 9'd4;
    parameter ap_ST_fsm_state4 = 9'd8;
    parameter ap_ST_fsm_state5 = 9'd16;
    parameter ap_ST_fsm_state6 = 9'd32;
    parameter ap_ST_fsm_state7 = 9'd64;
    parameter ap_ST_fsm_state8 = 9'd128;
    parameter ap_ST_fsm_state9 = 9'd256;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [62:0] in_val;
    input [11:0] prescale;
    output [63:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[63:0] ap_return;

    (* fsm_encoding = "none" *) reg   [8:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire    ap_CS_fsm_state3;
    wire   [14:0] trunc_ln408_fu_168_p1;
    reg   [14:0] trunc_ln408_reg_422;
    wire   [31:0] out_bits_3_fu_184_p3;
    reg   [31:0] out_bits_3_reg_436;
    wire    ap_CS_fsm_state5;
    wire   [0:0] icmp_ln433_fu_208_p2;
    reg   [0:0] icmp_ln433_reg_453;
    wire    ap_CS_fsm_state7;
    wire   [0:0] grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_return;
    reg   [0:0] targetBlock_reg_458;
    wire    ap_CS_fsm_state8;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_done;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_idle;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_ready;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out_ap_vld;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_done;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_idle;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_ready;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_2_2_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_2_2_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_1_2_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_1_2_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_0_21_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_0_21_out_ap_vld;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_done;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_idle;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_ready;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_2_05_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_2_05_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_1_04_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_1_04_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_0_03_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_0_03_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_3_02_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_3_02_out_ap_vld;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_done;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_idle;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_ready;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out_ap_vld;
    wire   [61:0] grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out_ap_vld;
    wire   [31:0] grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out_ap_vld;
    wire   [61:0] grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out;
    wire    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out_ap_vld;
    reg    grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg;
    reg   [31:0] out_bits_2_1_loc_fu_96;
    wire    ap_CS_fsm_state2;
    reg   [31:0] out_bits_1_1_loc_fu_92;
    reg   [31:0] out_bits_0_1_loc_fu_88;
    reg    grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg;
    wire    ap_CS_fsm_state4;
    reg    grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg;
    wire    ap_CS_fsm_state6;
    reg    grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg;
    reg   [31:0] shift_loc_fu_56;
    reg   [61:0] in_shift_loc_fu_52;
    reg   [31:0] shift_1_loc_fu_48;
    reg   [61:0] in_shift_1_loc_fu_44;
    wire    ap_CS_fsm_state9;
    wire   [11:0] sub_ln432_fu_232_p2;
    wire  signed [31:0] sext_ln432_fu_238_p1;
    wire   [31:0] select_ln421_fu_225_p3;
    wire   [31:0] newexp_fu_242_p2;
    wire   [0:0] tmp_fu_248_p3;
    wire   [51:0] tmp_19_fu_261_p4;
    wire   [51:0] tmp_20_fu_271_p4;
    wire   [0:0] or_ln433_fu_256_p2;
    wire   [51:0] select_ln421_1_fu_281_p3;
    wire   [10:0] empty_fu_288_p1;
    wire   [10:0] out_exp_fu_300_p3;
    wire   [51:0] significand_fu_292_p3;
    wire   [63:0] t_fu_308_p4;
    wire   [63:0] bitcast_ln497_fu_318_p1;
    reg   [63:0] ap_return_preg;
    reg   [8:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    reg    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    reg    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    reg    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    reg    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 9'd1;
        #0 grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg = 1'b0;
        #0 grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg = 1'b0;
        #0 grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg = 1'b0;
        #0 grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg = 1'b0;
        #0 ap_return_preg = 64'd0;
    end

    main_scaled_fixed2ieee_63_1_Pipeline_1 grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start),
        .ap_done(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_done),
        .ap_idle(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_idle),
        .ap_ready(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_ready),
        .out_bits_2_1_out(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out),
        .out_bits_2_1_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out_ap_vld),
        .out_bits_1_1_out(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out),
        .out_bits_1_1_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out_ap_vld),
        .out_bits_0_1_out(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out),
        .out_bits_0_1_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out_ap_vld)
    );

    main_scaled_fixed2ieee_63_1_Pipeline_2 grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start),
        .ap_done(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_done),
        .ap_idle(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_idle),
        .ap_ready(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_ready),
        .out_bits_2_1_reload(out_bits_2_1_loc_fu_96),
        .out_bits_1_1_reload(out_bits_1_1_loc_fu_92),
        .out_bits_0_1_reload(out_bits_0_1_loc_fu_88),
        .in_val(in_val),
        .out_bits_2_2_out(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_2_2_out),
        .out_bits_2_2_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_2_2_out_ap_vld),
        .out_bits_1_2_out(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_1_2_out),
        .out_bits_1_2_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_1_2_out_ap_vld),
        .out_bits_0_21_out(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_0_21_out),
        .out_bits_0_21_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_0_21_out_ap_vld)
    );

    main_scaled_fixed2ieee_63_1_Pipeline_3 grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start),
        .ap_done(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_done),
        .ap_idle(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_idle),
        .ap_ready(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_ready),
        .out_bits_0_21_reload(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_0_21_out),
        .out_bits_1_2_reload(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_1_2_out),
        .out_bits_2_2_reload(grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_out_bits_2_2_out),
        .out_bits_3(out_bits_3_reg_436),
        .c_2_05_out(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_2_05_out),
        .c_2_05_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_2_05_out_ap_vld),
        .c_1_04_out(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_1_04_out),
        .c_1_04_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_1_04_out_ap_vld),
        .c_0_03_out(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_0_03_out),
        .c_0_03_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_0_03_out_ap_vld),
        .c_3_02_out(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_3_02_out),
        .c_3_02_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_3_02_out_ap_vld)
    );

    main_scaled_fixed2ieee_63_1_Pipeline_4 grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start),
        .ap_done(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_done),
        .ap_idle(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_idle),
        .ap_ready(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_ready),
        .in_val(in_val),
        .c_0_03_reload(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_0_03_out),
        .c_1_04_reload(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_1_04_out),
        .c_2_05_reload(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_2_05_out),
        .c_3_02_reload(grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_c_3_02_out),
        .shift_out(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out),
        .shift_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out_ap_vld),
        .in_shift_out(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out),
        .in_shift_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out_ap_vld),
        .shift_1_out(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out),
        .shift_1_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out_ap_vld),
        .in_shift_1_out(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out),
        .in_shift_1_out_ap_vld(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out_ap_vld),
        .ap_return(grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_return)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg[0]  <= 1'b0;
            ap_return_preg[1]  <= 1'b0;
            ap_return_preg[2]  <= 1'b0;
            ap_return_preg[3]  <= 1'b0;
            ap_return_preg[4]  <= 1'b0;
            ap_return_preg[5]  <= 1'b0;
            ap_return_preg[6]  <= 1'b0;
            ap_return_preg[7]  <= 1'b0;
            ap_return_preg[8]  <= 1'b0;
            ap_return_preg[9]  <= 1'b0;
            ap_return_preg[10] <= 1'b0;
            ap_return_preg[11] <= 1'b0;
            ap_return_preg[12] <= 1'b0;
            ap_return_preg[13] <= 1'b0;
            ap_return_preg[14] <= 1'b0;
            ap_return_preg[15] <= 1'b0;
            ap_return_preg[16] <= 1'b0;
            ap_return_preg[17] <= 1'b0;
            ap_return_preg[18] <= 1'b0;
            ap_return_preg[19] <= 1'b0;
            ap_return_preg[20] <= 1'b0;
            ap_return_preg[21] <= 1'b0;
            ap_return_preg[22] <= 1'b0;
            ap_return_preg[23] <= 1'b0;
            ap_return_preg[24] <= 1'b0;
            ap_return_preg[25] <= 1'b0;
            ap_return_preg[26] <= 1'b0;
            ap_return_preg[27] <= 1'b0;
            ap_return_preg[28] <= 1'b0;
            ap_return_preg[29] <= 1'b0;
            ap_return_preg[30] <= 1'b0;
            ap_return_preg[31] <= 1'b0;
            ap_return_preg[32] <= 1'b0;
            ap_return_preg[33] <= 1'b0;
            ap_return_preg[34] <= 1'b0;
            ap_return_preg[35] <= 1'b0;
            ap_return_preg[36] <= 1'b0;
            ap_return_preg[37] <= 1'b0;
            ap_return_preg[38] <= 1'b0;
            ap_return_preg[39] <= 1'b0;
            ap_return_preg[40] <= 1'b0;
            ap_return_preg[41] <= 1'b0;
            ap_return_preg[42] <= 1'b0;
            ap_return_preg[43] <= 1'b0;
            ap_return_preg[44] <= 1'b0;
            ap_return_preg[45] <= 1'b0;
            ap_return_preg[46] <= 1'b0;
            ap_return_preg[47] <= 1'b0;
            ap_return_preg[48] <= 1'b0;
            ap_return_preg[49] <= 1'b0;
            ap_return_preg[50] <= 1'b0;
            ap_return_preg[51] <= 1'b0;
            ap_return_preg[52] <= 1'b0;
            ap_return_preg[53] <= 1'b0;
            ap_return_preg[54] <= 1'b0;
            ap_return_preg[55] <= 1'b0;
            ap_return_preg[56] <= 1'b0;
            ap_return_preg[57] <= 1'b0;
            ap_return_preg[58] <= 1'b0;
            ap_return_preg[59] <= 1'b0;
            ap_return_preg[60] <= 1'b0;
            ap_return_preg[61] <= 1'b0;
            ap_return_preg[62] <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state9)) begin
                ap_return_preg[62 : 0] <= bitcast_ln497_fu_318_p1[62 : 0];
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg <= 1'b1;
            end else if ((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_ready == 1'b1)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg <= 1'b1;
            end else if ((grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_ready == 1'b1)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state5)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg <= 1'b1;
            end else if ((grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_ready == 1'b1)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state7)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg <= 1'b1;
            end else if ((grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_ready == 1'b1)) begin
                grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state7)) begin
            icmp_ln433_reg_453 <= icmp_ln433_fu_208_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out_ap_vld == 1'b1))) begin
            in_shift_1_loc_fu_44 <= grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out_ap_vld == 1'b1))) begin
            in_shift_loc_fu_52 <= grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_in_shift_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
            out_bits_0_1_loc_fu_88 <= grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_0_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
            out_bits_1_1_loc_fu_92 <= grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_1_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
            out_bits_2_1_loc_fu_96 <= grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_out_bits_2_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state5)) begin
            out_bits_3_reg_436[31 : 17] <= out_bits_3_fu_184_p3[31 : 17];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out_ap_vld == 1'b1))) begin
            shift_1_loc_fu_48 <= grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_1_out;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_state8) & (grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out_ap_vld == 1'b1))) begin
            shift_loc_fu_56 <= grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_shift_out;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            targetBlock_reg_458 <= grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_return;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            trunc_ln408_reg_422 <= trunc_ln408_fu_168_p1;
        end
    end

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_done == 1'b0)) begin
            ap_ST_fsm_state2_blk = 1'b1;
        end else begin
            ap_ST_fsm_state2_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state3_blk = 1'b0;

    always @(*) begin
        if ((grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_done == 1'b0)) begin
            ap_ST_fsm_state4_blk = 1'b1;
        end else begin
            ap_ST_fsm_state4_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state5_blk = 1'b0;

    always @(*) begin
        if ((grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_done == 1'b0)) begin
            ap_ST_fsm_state6_blk = 1'b1;
        end else begin
            ap_ST_fsm_state6_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state7_blk = 1'b0;

    always @(*) begin
        if ((grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_done == 1'b0)) begin
            ap_ST_fsm_state8_blk = 1'b1;
        end else begin
            ap_ST_fsm_state8_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state9_blk = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state9) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_return = bitcast_ln497_fu_318_p1;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                if (((grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                if (((grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state4))) begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                if (((grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state6))) begin
                    ap_NS_fsm = ap_ST_fsm_state7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state6;
                end
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                if (((1'b1 == ap_CS_fsm_state8) & (grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_done == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state8;
                end
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign bitcast_ln497_fu_318_p1 = t_fu_308_p4;

    assign empty_fu_288_p1 = newexp_fu_242_p2[10:0];

    assign grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start = grp_scaled_fixed2ieee_63_1_Pipeline_1_fu_112_ap_start_reg;

    assign grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start = grp_scaled_fixed2ieee_63_1_Pipeline_2_fu_119_ap_start_reg;

    assign grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start = grp_scaled_fixed2ieee_63_1_Pipeline_3_fu_131_ap_start_reg;

    assign grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start = grp_scaled_fixed2ieee_63_1_Pipeline_4_fu_143_ap_start_reg;

    assign icmp_ln433_fu_208_p2 = ((in_val == 63'd0) ? 1'b1 : 1'b0);

    assign newexp_fu_242_p2 = ($signed(sext_ln432_fu_238_p1) - $signed(select_ln421_fu_225_p3));

    assign or_ln433_fu_256_p2 = (tmp_fu_248_p3 | icmp_ln433_reg_453);

    assign out_bits_3_fu_184_p3 = {{trunc_ln408_reg_422}, {17'd65536}};

    assign out_exp_fu_300_p3 = ((or_ln433_fu_256_p2[0:0] == 1'b1) ? 11'd0 : empty_fu_288_p1);

    assign select_ln421_1_fu_281_p3 = ((targetBlock_reg_458[0:0] == 1'b1) ? tmp_19_fu_261_p4 : tmp_20_fu_271_p4);

    assign select_ln421_fu_225_p3 = ((targetBlock_reg_458[0:0] == 1'b1) ? shift_loc_fu_56 : shift_1_loc_fu_48);

    assign sext_ln432_fu_238_p1 = $signed(sub_ln432_fu_232_p2);

    assign significand_fu_292_p3 = ((or_ln433_fu_256_p2[0:0] == 1'b1) ? 52'd0 : select_ln421_1_fu_281_p3);

    assign sub_ln432_fu_232_p2 = (12'd1023 - prescale);

    assign t_fu_308_p4 = {{{{1'd0}, {out_exp_fu_300_p3}}}, {significand_fu_292_p3}};

    assign tmp_19_fu_261_p4 = {{in_shift_loc_fu_52[61:10]}};

    assign tmp_20_fu_271_p4 = {{in_shift_1_loc_fu_44[61:10]}};

    assign tmp_fu_248_p3 = newexp_fu_242_p2[32'd31];

    assign trunc_ln408_fu_168_p1 = in_val[14:0];

    always @(posedge ap_clk) begin
        out_bits_3_reg_436[16:0] <= 17'b10000000000000000;
        ap_return_preg[63] <= 1'b0;
    end

endmodule  //main_scaled_fixed2ieee_63_1_s
