/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_42_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    sum_out,
    sum_out_ap_vld
);

    parameter ap_ST_fsm_pp0_stage0 = 7'd1;
    parameter ap_ST_fsm_pp0_stage1 = 7'd2;
    parameter ap_ST_fsm_pp0_stage2 = 7'd4;
    parameter ap_ST_fsm_pp0_stage3 = 7'd8;
    parameter ap_ST_fsm_pp0_stage4 = 7'd16;
    parameter ap_ST_fsm_pp0_stage5 = 7'd32;
    parameter ap_ST_fsm_pp0_stage6 = 7'd64;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [63:0] sum_out;
    output sum_out_ap_vld;

    reg ap_idle;
    reg sum_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [6:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_subdone;
    reg   [0:0] icmp_ln42_reg_182;
    reg    ap_condition_exit_pp0_iter0_stage6;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    wire   [0:0] icmp_ln42_fu_103_p2;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter1_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter2_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter3_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter4_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter5_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter6_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter7_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter8_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter9_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter10_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter11_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter12_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter13_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter14_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter15_reg;
    reg   [0:0] icmp_ln42_reg_182_pp0_iter16_reg;
    wire   [63:0] grp_fu_77_p1;
    reg   [63:0] conv_reg_191;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire   [63:0] grp_fu_72_p2;
    reg   [63:0] actual_value_reg_196;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    reg   [63:0] actual_value_reg_196_pp0_iter10_reg;
    wire   [63:0] grp_fu_61_p2;
    reg   [63:0] setpoint_reg_202;
    reg   [63:0] error_reg_207;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [63:0] error_reg_207_pp0_iter12_reg;
    reg   [63:0] error_reg_207_pp0_iter13_reg;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    reg   [63:0] controller_integral_1_reg_224;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    reg   [63:0] derivative_reg_230;
    wire   [63:0] grp_fu_66_p2;
    reg   [63:0] mul4_i_reg_235;
    reg   [63:0] mul6_i_reg_240;
    reg   [63:0] mul6_i_reg_240_pp0_iter14_reg;
    reg   [63:0] add5_i_reg_245;
    reg   [63:0] output_reg_250;
    wire    ap_block_pp0_stage6_11001;
    reg   [63:0] sum_1_reg_260;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage1_subdone;
    reg   [63:0] sum_fu_38;
    reg   [63:0] ap_sig_allocacmp_sum_load;
    wire    ap_block_pp0_stage1;
    wire    ap_loop_init;
    reg   [9:0] i_fu_42;
    wire   [9:0] i_2_fu_109_p2;
    reg   [9:0] ap_sig_allocacmp_i_1;
    wire    ap_block_pp0_stage0;
    reg   [63:0] controller_integral_fu_46;
    reg   [63:0] ap_sig_allocacmp_controller_integral_load;
    wire    ap_block_pp0_stage4;
    reg   [63:0] controller_previous_error_fu_50;
    wire    ap_block_pp0_stage5;
    wire    ap_block_pp0_stage1_01001;
    reg   [63:0] grp_fu_61_p0;
    reg   [63:0] grp_fu_61_p1;
    wire    ap_block_pp0_stage2;
    wire    ap_block_pp0_stage3;
    wire    ap_block_pp0_stage6;
    reg   [63:0] grp_fu_66_p0;
    reg   [63:0] grp_fu_66_p1;
    wire   [31:0] grp_fu_77_p0;
    reg   [1:0] grp_fu_61_opcode;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage6_00001;
    wire    ap_block_pp0_stage0_00001;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage5_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    reg    ap_condition_exit_pp0_iter16_stage1;
    reg    ap_idle_pp0_0to15;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg    ap_loop_exit_ready_pp0_iter10_reg;
    reg    ap_loop_exit_ready_pp0_iter11_reg;
    reg    ap_loop_exit_ready_pp0_iter12_reg;
    reg    ap_loop_exit_ready_pp0_iter13_reg;
    reg    ap_loop_exit_ready_pp0_iter14_reg;
    reg    ap_loop_exit_ready_pp0_iter15_reg;
    reg    ap_loop_exit_ready_pp0_iter16_reg;
    reg   [6:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to17;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 7'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 sum_fu_38 = 64'd0;
        #0 i_fu_42 = 10'd0;
        #0 controller_integral_fu_46 = 64'd0;
        #0 controller_previous_error_fu_50 = 64'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_dadddsub_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_U1 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_61_p0),
        .din1(grp_fu_61_p1),
        .opcode(grp_fu_61_opcode),
        .ce(1'b1),
        .dout(grp_fu_61_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U2 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_66_p0),
        .din1(grp_fu_66_p1),
        .ce(1'b1),
        .dout(grp_fu_66_p2)
    );

    main_ddiv_64ns_64ns_64_59_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(59),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) ddiv_64ns_64ns_64_59_no_dsp_1_U3 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(conv_reg_191),
        .din1(64'd4621819117588971520),
        .ce(1'b1),
        .dout(grp_fu_72_p2)
    );

    main_sitodp_32ns_64_6_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(6),
        .din0_WIDTH(32),
        .dout_WIDTH(64)
    ) sitodp_32ns_64_6_no_dsp_1_U4 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_77_p0),
        .ce(1'b1),
        .dout(grp_fu_77_p1)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage6),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_loop_exit_ready_pp0_iter16_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage6)) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                ap_enable_reg_pp0_iter17 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage6_subdone) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter13_reg <= ap_loop_exit_ready_pp0_iter12_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter14_reg <= ap_loop_exit_ready_pp0_iter13_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter15_reg <= ap_loop_exit_ready_pp0_iter14_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter16_reg <= ap_loop_exit_ready_pp0_iter15_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage6_11001) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            controller_integral_fu_46 <= 64'd0;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            controller_integral_fu_46 <= controller_integral_1_reg_224;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            controller_previous_error_fu_50 <= 64'd0;
        end else if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            controller_previous_error_fu_50 <= error_reg_207;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln42_fu_103_p2 == 1'd0))) begin
                i_fu_42 <= i_2_fu_109_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                i_fu_42 <= 10'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            sum_fu_38 <= 64'd0;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            sum_fu_38 <= sum_1_reg_260;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            actual_value_reg_196 <= grp_fu_72_p2;
            actual_value_reg_196_pp0_iter10_reg <= actual_value_reg_196;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            add5_i_reg_245 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            controller_integral_1_reg_224 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage5_11001) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            conv_reg_191 <= grp_fu_77_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            derivative_reg_230 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            error_reg_207 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            error_reg_207_pp0_iter12_reg <= error_reg_207;
            error_reg_207_pp0_iter13_reg <= error_reg_207_pp0_iter12_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            icmp_ln42_reg_182 <= icmp_ln42_fu_103_p2;
            icmp_ln42_reg_182_pp0_iter10_reg <= icmp_ln42_reg_182_pp0_iter9_reg;
            icmp_ln42_reg_182_pp0_iter11_reg <= icmp_ln42_reg_182_pp0_iter10_reg;
            icmp_ln42_reg_182_pp0_iter12_reg <= icmp_ln42_reg_182_pp0_iter11_reg;
            icmp_ln42_reg_182_pp0_iter13_reg <= icmp_ln42_reg_182_pp0_iter12_reg;
            icmp_ln42_reg_182_pp0_iter14_reg <= icmp_ln42_reg_182_pp0_iter13_reg;
            icmp_ln42_reg_182_pp0_iter15_reg <= icmp_ln42_reg_182_pp0_iter14_reg;
            icmp_ln42_reg_182_pp0_iter16_reg <= icmp_ln42_reg_182_pp0_iter15_reg;
            icmp_ln42_reg_182_pp0_iter1_reg <= icmp_ln42_reg_182;
            icmp_ln42_reg_182_pp0_iter2_reg <= icmp_ln42_reg_182_pp0_iter1_reg;
            icmp_ln42_reg_182_pp0_iter3_reg <= icmp_ln42_reg_182_pp0_iter2_reg;
            icmp_ln42_reg_182_pp0_iter4_reg <= icmp_ln42_reg_182_pp0_iter3_reg;
            icmp_ln42_reg_182_pp0_iter5_reg <= icmp_ln42_reg_182_pp0_iter4_reg;
            icmp_ln42_reg_182_pp0_iter6_reg <= icmp_ln42_reg_182_pp0_iter5_reg;
            icmp_ln42_reg_182_pp0_iter7_reg <= icmp_ln42_reg_182_pp0_iter6_reg;
            icmp_ln42_reg_182_pp0_iter8_reg <= icmp_ln42_reg_182_pp0_iter7_reg;
            icmp_ln42_reg_182_pp0_iter9_reg <= icmp_ln42_reg_182_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            mul4_i_reg_235 <= grp_fu_66_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul6_i_reg_240 <= grp_fu_66_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            mul6_i_reg_240_pp0_iter14_reg <= mul6_i_reg_240;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            output_reg_250 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            setpoint_reg_202 <= grp_fu_61_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            sum_1_reg_260 <= grp_fu_61_p2;
        end
    end

    always @(*) begin
        if (((icmp_ln42_reg_182 == 1'd1) & (1'b0 == ap_block_pp0_stage6_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_condition_exit_pp0_iter0_stage6 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage6 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln42_reg_182_pp0_iter16_reg == 1'd1))) begin
            ap_condition_exit_pp0_iter16_stage1 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter16_stage1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_loop_exit_ready_pp0_iter16_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to15 = 1'b1;
        end else begin
            ap_idle_pp0_0to15 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to17 = 1'b1;
        end else begin
            ap_idle_pp0_1to17 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage6_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            ap_sig_allocacmp_controller_integral_load = controller_integral_1_reg_224;
        end else begin
            ap_sig_allocacmp_controller_integral_load = controller_integral_fu_46;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_sig_allocacmp_i_1 = 10'd0;
        end else begin
            ap_sig_allocacmp_i_1 = i_fu_42;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter17 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_sig_allocacmp_sum_load = sum_1_reg_260;
        end else begin
            ap_sig_allocacmp_sum_load = sum_fu_38;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_61_opcode = 2'd1;
        end else if ((((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_61_opcode = 2'd0;
        end else begin
            grp_fu_61_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_61_p0 = ap_sig_allocacmp_sum_load;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_61_p0 = add5_i_reg_245;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_61_p0 = error_reg_207_pp0_iter13_reg;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_61_p0 = error_reg_207;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_61_p0 = ap_sig_allocacmp_controller_integral_load;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_61_p0 = setpoint_reg_202;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_61_p0 = actual_value_reg_196;
        end else begin
            grp_fu_61_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter16 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_61_p1 = output_reg_250;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter15 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            grp_fu_61_p1 = mul6_i_reg_240_pp0_iter14_reg;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter13 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            grp_fu_61_p1 = mul4_i_reg_235;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_61_p1 = controller_previous_error_fu_50;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter11 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_61_p1 = error_reg_207;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter10 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_61_p1 = actual_value_reg_196_pp0_iter10_reg;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_61_p1 = 64'd4607182418800017408;
        end else begin
            grp_fu_61_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter12 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                grp_fu_66_p0 = derivative_reg_230;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                grp_fu_66_p0 = controller_integral_1_reg_224;
            end else begin
                grp_fu_66_p0 = 'bx;
            end
        end else begin
            grp_fu_66_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter12 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                grp_fu_66_p1 = 64'd4576918229304087675;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                grp_fu_66_p1 = 64'd4591870180066957722;
            end else begin
                grp_fu_66_p1 = 'bx;
            end
        end else begin
            grp_fu_66_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln42_reg_182_pp0_iter16_reg == 1'd1))) begin
            sum_out_ap_vld = 1'b1;
        end else begin
            sum_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to17 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if (((ap_idle_pp0_0to15 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter16_stage1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage6;

    assign grp_fu_77_p0 = ap_sig_allocacmp_i_1;

    assign i_2_fu_109_p2 = (ap_sig_allocacmp_i_1 + 10'd1);

    assign icmp_ln42_fu_103_p2 = ((ap_sig_allocacmp_i_1 == 10'd1000) ? 1'b1 : 1'b0);

    assign sum_out = sum_fu_38;

endmodule  //main_main_Pipeline_VITIS_LOOP_42_1
