/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_atan2_generic_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    y_in,
    x_in,
    ap_return
);

    parameter ap_ST_fsm_state1 = 116'd1;
    parameter ap_ST_fsm_state2 = 116'd2;
    parameter ap_ST_fsm_state3 = 116'd4;
    parameter ap_ST_fsm_state4 = 116'd8;
    parameter ap_ST_fsm_state5 = 116'd16;
    parameter ap_ST_fsm_state6 = 116'd32;
    parameter ap_ST_fsm_state7 = 116'd64;
    parameter ap_ST_fsm_state8 = 116'd128;
    parameter ap_ST_fsm_state9 = 116'd256;
    parameter ap_ST_fsm_state10 = 116'd512;
    parameter ap_ST_fsm_state11 = 116'd1024;
    parameter ap_ST_fsm_state12 = 116'd2048;
    parameter ap_ST_fsm_state13 = 116'd4096;
    parameter ap_ST_fsm_state14 = 116'd8192;
    parameter ap_ST_fsm_state15 = 116'd16384;
    parameter ap_ST_fsm_state16 = 116'd32768;
    parameter ap_ST_fsm_state17 = 116'd65536;
    parameter ap_ST_fsm_state18 = 116'd131072;
    parameter ap_ST_fsm_state19 = 116'd262144;
    parameter ap_ST_fsm_state20 = 116'd524288;
    parameter ap_ST_fsm_state21 = 116'd1048576;
    parameter ap_ST_fsm_state22 = 116'd2097152;
    parameter ap_ST_fsm_state23 = 116'd4194304;
    parameter ap_ST_fsm_state24 = 116'd8388608;
    parameter ap_ST_fsm_state25 = 116'd16777216;
    parameter ap_ST_fsm_state26 = 116'd33554432;
    parameter ap_ST_fsm_state27 = 116'd67108864;
    parameter ap_ST_fsm_state28 = 116'd134217728;
    parameter ap_ST_fsm_state29 = 116'd268435456;
    parameter ap_ST_fsm_state30 = 116'd536870912;
    parameter ap_ST_fsm_state31 = 116'd1073741824;
    parameter ap_ST_fsm_state32 = 116'd2147483648;
    parameter ap_ST_fsm_state33 = 116'd4294967296;
    parameter ap_ST_fsm_state34 = 116'd8589934592;
    parameter ap_ST_fsm_state35 = 116'd17179869184;
    parameter ap_ST_fsm_state36 = 116'd34359738368;
    parameter ap_ST_fsm_state37 = 116'd68719476736;
    parameter ap_ST_fsm_state38 = 116'd137438953472;
    parameter ap_ST_fsm_state39 = 116'd274877906944;
    parameter ap_ST_fsm_state40 = 116'd549755813888;
    parameter ap_ST_fsm_state41 = 116'd1099511627776;
    parameter ap_ST_fsm_state42 = 116'd2199023255552;
    parameter ap_ST_fsm_state43 = 116'd4398046511104;
    parameter ap_ST_fsm_state44 = 116'd8796093022208;
    parameter ap_ST_fsm_state45 = 116'd17592186044416;
    parameter ap_ST_fsm_state46 = 116'd35184372088832;
    parameter ap_ST_fsm_state47 = 116'd70368744177664;
    parameter ap_ST_fsm_state48 = 116'd140737488355328;
    parameter ap_ST_fsm_state49 = 116'd281474976710656;
    parameter ap_ST_fsm_state50 = 116'd562949953421312;
    parameter ap_ST_fsm_state51 = 116'd1125899906842624;
    parameter ap_ST_fsm_state52 = 116'd2251799813685248;
    parameter ap_ST_fsm_state53 = 116'd4503599627370496;
    parameter ap_ST_fsm_state54 = 116'd9007199254740992;
    parameter ap_ST_fsm_state55 = 116'd18014398509481984;
    parameter ap_ST_fsm_state56 = 116'd36028797018963968;
    parameter ap_ST_fsm_state57 = 116'd72057594037927936;
    parameter ap_ST_fsm_state58 = 116'd144115188075855872;
    parameter ap_ST_fsm_state59 = 116'd288230376151711744;
    parameter ap_ST_fsm_state60 = 116'd576460752303423488;
    parameter ap_ST_fsm_state61 = 116'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 116'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 116'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 116'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 116'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 116'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 116'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 116'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 116'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 116'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 116'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 116'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 116'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 116'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 116'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 116'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 116'd75557863725914323419136;
    parameter ap_ST_fsm_state78 = 116'd151115727451828646838272;
    parameter ap_ST_fsm_state79 = 116'd302231454903657293676544;
    parameter ap_ST_fsm_state80 = 116'd604462909807314587353088;
    parameter ap_ST_fsm_state81 = 116'd1208925819614629174706176;
    parameter ap_ST_fsm_state82 = 116'd2417851639229258349412352;
    parameter ap_ST_fsm_state83 = 116'd4835703278458516698824704;
    parameter ap_ST_fsm_state84 = 116'd9671406556917033397649408;
    parameter ap_ST_fsm_state85 = 116'd19342813113834066795298816;
    parameter ap_ST_fsm_state86 = 116'd38685626227668133590597632;
    parameter ap_ST_fsm_state87 = 116'd77371252455336267181195264;
    parameter ap_ST_fsm_state88 = 116'd154742504910672534362390528;
    parameter ap_ST_fsm_state89 = 116'd309485009821345068724781056;
    parameter ap_ST_fsm_state90 = 116'd618970019642690137449562112;
    parameter ap_ST_fsm_state91 = 116'd1237940039285380274899124224;
    parameter ap_ST_fsm_state92 = 116'd2475880078570760549798248448;
    parameter ap_ST_fsm_state93 = 116'd4951760157141521099596496896;
    parameter ap_ST_fsm_state94 = 116'd9903520314283042199192993792;
    parameter ap_ST_fsm_state95 = 116'd19807040628566084398385987584;
    parameter ap_ST_fsm_state96 = 116'd39614081257132168796771975168;
    parameter ap_ST_fsm_state97 = 116'd79228162514264337593543950336;
    parameter ap_ST_fsm_state98 = 116'd158456325028528675187087900672;
    parameter ap_ST_fsm_state99 = 116'd316912650057057350374175801344;
    parameter ap_ST_fsm_state100 = 116'd633825300114114700748351602688;
    parameter ap_ST_fsm_state101 = 116'd1267650600228229401496703205376;
    parameter ap_ST_fsm_state102 = 116'd2535301200456458802993406410752;
    parameter ap_ST_fsm_state103 = 116'd5070602400912917605986812821504;
    parameter ap_ST_fsm_state104 = 116'd10141204801825835211973625643008;
    parameter ap_ST_fsm_state105 = 116'd20282409603651670423947251286016;
    parameter ap_ST_fsm_state106 = 116'd40564819207303340847894502572032;
    parameter ap_ST_fsm_state107 = 116'd81129638414606681695789005144064;
    parameter ap_ST_fsm_state108 = 116'd162259276829213363391578010288128;
    parameter ap_ST_fsm_state109 = 116'd324518553658426726783156020576256;
    parameter ap_ST_fsm_state110 = 116'd649037107316853453566312041152512;
    parameter ap_ST_fsm_state111 = 116'd1298074214633706907132624082305024;
    parameter ap_ST_fsm_state112 = 116'd2596148429267413814265248164610048;
    parameter ap_ST_fsm_state113 = 116'd5192296858534827628530496329220096;
    parameter ap_ST_fsm_state114 = 116'd10384593717069655257060992658440192;
    parameter ap_ST_fsm_state115 = 116'd20769187434139310514121985316880384;
    parameter ap_ST_fsm_state116 = 116'd41538374868278621028243970633760768;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] y_in;
    input [63:0] x_in;
    output [63:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[63:0] ap_return;

    (* fsm_encoding = "none" *) reg   [115:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire   [0:0] icmp_ln655_fu_186_p2;
    reg   [0:0] icmp_ln655_reg_618;
    wire   [51:0] trunc_ln505_fu_208_p1;
    reg   [51:0] trunc_ln505_reg_625;
    wire   [51:0] trunc_ln505_2_fu_212_p1;
    reg   [51:0] trunc_ln505_2_reg_630;
    wire   [0:0] tmp_fu_216_p3;
    reg   [0:0] tmp_reg_635;
    wire   [10:0] select_ln695_fu_230_p3;
    reg   [10:0] select_ln695_reg_640;
    wire   [88:0] y_3_fu_266_p3;
    reg   [88:0] y_3_reg_645;
    wire    ap_CS_fsm_state2;
    wire   [85:0] x_fu_273_p4;
    reg   [85:0] x_reg_650;
    wire    ap_CS_fsm_state3;
    wire   [0:0] tmp_28_fu_292_p3;
    reg   [0:0] tmp_28_reg_658;
    wire    ap_CS_fsm_state53;
    wire   [85:0] select_ln702_fu_306_p3;
    reg   [85:0] select_ln702_reg_663;
    reg   [63:0] tmp_s_reg_671;
    wire   [21:0] trunc_ln702_1_fu_324_p1;
    reg   [21:0] trunc_ln702_1_reg_677;
    wire   [10:0] trunc_ln702_3_fu_377_p1;
    reg   [10:0] trunc_ln702_3_reg_682;
    wire    ap_CS_fsm_state54;
    wire   [31:0] sub_ln702_1_fu_381_p2;
    reg   [31:0] sub_ln702_1_reg_687;
    wire   [6:0] trunc_ln702_4_fu_387_p1;
    reg   [6:0] trunc_ln702_4_reg_694;
    wire   [85:0] lshr_ln702_2_fu_400_p2;
    reg   [85:0] lshr_ln702_2_reg_699;
    wire    ap_CS_fsm_state55;
    wire   [1:0] or_ln_fu_476_p3;
    reg   [1:0] or_ln_reg_704;
    wire    ap_CS_fsm_state56;
    wire   [0:0] icmp_ln702_4_fu_484_p2;
    reg   [0:0] icmp_ln702_4_reg_709;
    wire   [85:0] lshr_ln702_fu_499_p2;
    reg   [85:0] lshr_ln702_reg_714;
    wire   [85:0] shl_ln702_fu_513_p2;
    reg   [85:0] shl_ln702_reg_719;
    reg   [62:0] lshr_ln702_1_reg_724;
    wire    ap_CS_fsm_state57;
    reg   [0:0] tmp_31_reg_729;
    wire   [63:0] bitcast_ln753_fu_598_p1;
    wire    ap_CS_fsm_state58;
    wire    grp_atan2_generic_double_Pipeline_1_fu_128_ap_start;
    wire    grp_atan2_generic_double_Pipeline_1_fu_128_ap_done;
    wire    grp_atan2_generic_double_Pipeline_1_fu_128_ap_idle;
    wire    grp_atan2_generic_double_Pipeline_1_fu_128_ap_ready;
    wire   [85:0] grp_atan2_generic_double_Pipeline_1_fu_128_z_out;
    wire    grp_atan2_generic_double_Pipeline_1_fu_128_z_out_ap_vld;
    wire   [63:0] grp_fu_137_p2;
    reg   [63:0] ap_phi_mux_retval_0_phi_fu_116_p8;
    reg   [63:0] retval_0_reg_112;
    wire    ap_CS_fsm_state116;
    wire   [0:0] icmp_ln662_fu_192_p2;
    wire   [0:0] icmp_ln702_fu_286_p2;
    reg    grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg;
    wire    ap_CS_fsm_state4;
    wire   [63:0] data_fu_144_p1;
    wire   [63:0] data_5_fu_158_p1;
    wire   [10:0] fps_y_exp_fu_162_p4;
    wire   [11:0] zext_ln655_fu_172_p1;
    wire   [10:0] fps_x_exp_fu_148_p4;
    wire   [11:0] add_ln655_fu_176_p2;
    wire   [11:0] zext_ln655_1_fu_182_p1;
    wire   [11:0] d_exp_fu_198_p2;
    wire   [10:0] trunc_ln688_fu_204_p1;
    wire   [10:0] sub_ln695_fu_224_p2;
    wire   [85:0] y_fu_238_p4;
    wire   [88:0] zext_ln681_fu_247_p1;
    wire   [88:0] zext_ln695_fu_251_p1;
    wire   [88:0] shl_ln695_fu_254_p2;
    wire   [88:0] lshr_ln695_fu_260_p2;
    wire   [85:0] sub_ln702_fu_300_p2;
    reg   [63:0] tmp_12_fu_328_p3;
    wire   [63:0] tmp_14_fu_344_p3;
    reg   [63:0] tmp_15_fu_351_p3;
    wire   [31:0] trunc_ln702_2_fu_359_p1;
    wire   [31:0] trunc_ln702_fu_335_p1;
    wire   [0:0] icmp_ln702_1_fu_339_p2;
    wire   [31:0] add_ln702_fu_363_p2;
    wire   [31:0] select_ln702_1_fu_369_p3;
    wire   [6:0] sub_ln702_4_fu_391_p2;
    wire   [85:0] zext_ln702_4_fu_396_p1;
    wire   [31:0] add_ln702_1_fu_406_p2;
    wire   [30:0] tmp_29_fu_411_p4;
    wire   [85:0] and_ln702_2_fu_427_p2;
    wire   [0:0] icmp_ln702_2_fu_421_p2;
    wire   [0:0] icmp_ln702_3_fu_431_p2;
    wire   [0:0] tmp_30_fu_443_p3;
    wire   [0:0] bit_select27_i_i_fu_457_p3;
    wire   [0:0] xor_ln702_fu_451_p2;
    wire   [0:0] and_ln702_1_fu_464_p2;
    wire   [0:0] and_ln702_fu_437_p2;
    wire   [0:0] or_ln702_fu_470_p2;
    wire   [31:0] add_ln702_2_fu_490_p2;
    wire   [85:0] zext_ln702_fu_495_p1;
    wire   [31:0] sub_ln702_2_fu_504_p2;
    wire   [85:0] zext_ln702_1_fu_509_p1;
    wire   [63:0] trunc_ln702_5_fu_518_p1;
    wire   [63:0] trunc_ln702_6_fu_521_p1;
    wire   [63:0] select_ln702_2_fu_524_p3;
    wire   [63:0] zext_ln702_2_fu_531_p1;
    wire   [63:0] add_ln702_3_fu_534_p2;
    wire   [10:0] sub_ln702_3_fu_568_p2;
    wire   [10:0] select_ln702_3_fu_561_p3;
    wire   [10:0] add_ln702_4_fu_573_p2;
    wire   [63:0] zext_ln702_3_fu_558_p1;
    wire   [11:0] tmp_17_fu_579_p3;
    wire   [63:0] LD_fu_586_p5;
    reg   [63:0] ap_return_preg;
    reg   [115:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    reg    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_ST_fsm_state62_blk;
    wire    ap_ST_fsm_state63_blk;
    wire    ap_ST_fsm_state64_blk;
    wire    ap_ST_fsm_state65_blk;
    wire    ap_ST_fsm_state66_blk;
    wire    ap_ST_fsm_state67_blk;
    wire    ap_ST_fsm_state68_blk;
    wire    ap_ST_fsm_state69_blk;
    wire    ap_ST_fsm_state70_blk;
    wire    ap_ST_fsm_state71_blk;
    wire    ap_ST_fsm_state72_blk;
    wire    ap_ST_fsm_state73_blk;
    wire    ap_ST_fsm_state74_blk;
    wire    ap_ST_fsm_state75_blk;
    wire    ap_ST_fsm_state76_blk;
    wire    ap_ST_fsm_state77_blk;
    wire    ap_ST_fsm_state78_blk;
    wire    ap_ST_fsm_state79_blk;
    wire    ap_ST_fsm_state80_blk;
    wire    ap_ST_fsm_state81_blk;
    wire    ap_ST_fsm_state82_blk;
    wire    ap_ST_fsm_state83_blk;
    wire    ap_ST_fsm_state84_blk;
    wire    ap_ST_fsm_state85_blk;
    wire    ap_ST_fsm_state86_blk;
    wire    ap_ST_fsm_state87_blk;
    wire    ap_ST_fsm_state88_blk;
    wire    ap_ST_fsm_state89_blk;
    wire    ap_ST_fsm_state90_blk;
    wire    ap_ST_fsm_state91_blk;
    wire    ap_ST_fsm_state92_blk;
    wire    ap_ST_fsm_state93_blk;
    wire    ap_ST_fsm_state94_blk;
    wire    ap_ST_fsm_state95_blk;
    wire    ap_ST_fsm_state96_blk;
    wire    ap_ST_fsm_state97_blk;
    wire    ap_ST_fsm_state98_blk;
    wire    ap_ST_fsm_state99_blk;
    wire    ap_ST_fsm_state100_blk;
    wire    ap_ST_fsm_state101_blk;
    wire    ap_ST_fsm_state102_blk;
    wire    ap_ST_fsm_state103_blk;
    wire    ap_ST_fsm_state104_blk;
    wire    ap_ST_fsm_state105_blk;
    wire    ap_ST_fsm_state106_blk;
    wire    ap_ST_fsm_state107_blk;
    wire    ap_ST_fsm_state108_blk;
    wire    ap_ST_fsm_state109_blk;
    wire    ap_ST_fsm_state110_blk;
    wire    ap_ST_fsm_state111_blk;
    wire    ap_ST_fsm_state112_blk;
    wire    ap_ST_fsm_state113_blk;
    wire    ap_ST_fsm_state114_blk;
    wire    ap_ST_fsm_state115_blk;
    wire    ap_ST_fsm_state116_blk;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 116'd1;
        #0 grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg = 1'b0;
        #0 ap_return_preg = 64'd0;
    end

    main_atan2_generic_double_Pipeline_1 grp_atan2_generic_double_Pipeline_1_fu_128 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_atan2_generic_double_Pipeline_1_fu_128_ap_start),
        .ap_done(grp_atan2_generic_double_Pipeline_1_fu_128_ap_done),
        .ap_idle(grp_atan2_generic_double_Pipeline_1_fu_128_ap_idle),
        .ap_ready(grp_atan2_generic_double_Pipeline_1_fu_128_ap_ready),
        .y_1(y_3_reg_645),
        .zext_ln681(x_reg_650),
        .z_out(grp_atan2_generic_double_Pipeline_1_fu_128_z_out),
        .z_out_ap_vld(grp_atan2_generic_double_Pipeline_1_fu_128_z_out_ap_vld)
    );

    main_ddiv_64ns_64ns_64_59_no_dsp_1 #(
        .ID(1),
        .NUM_STAGE(59),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) ddiv_64ns_64ns_64_59_no_dsp_1_U15 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(y_in),
        .din1(x_in),
        .ce(1'b1),
        .dout(grp_fu_137_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_return_preg <= 64'd0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state116)) begin
                ap_return_preg <= ap_phi_mux_retval_0_phi_fu_116_p8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg <= 1'b1;
            end else if ((grp_atan2_generic_double_Pipeline_1_fu_128_ap_ready == 1'b1)) begin
                grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((((icmp_ln702_fu_286_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state53)) | ((icmp_ln662_fu_192_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1) & (icmp_ln655_fu_186_p2 == 1'd0) & (ap_start == 1'b1)))) begin
            retval_0_reg_112 <= 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state58)) begin
            retval_0_reg_112 <= bitcast_ln753_fu_598_p1;
        end else if (((1'b1 == ap_CS_fsm_state116) & (icmp_ln655_reg_618 == 1'd1))) begin
            retval_0_reg_112 <= grp_fu_137_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            icmp_ln655_reg_618 <= icmp_ln655_fu_186_p2;
            select_ln695_reg_640 <= select_ln695_fu_230_p3;
            tmp_reg_635 <= d_exp_fu_198_p2[32'd11];
            trunc_ln505_2_reg_630 <= trunc_ln505_2_fu_212_p1;
            trunc_ln505_reg_625 <= trunc_ln505_fu_208_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state56)) begin
            icmp_ln702_4_reg_709 <= icmp_ln702_4_fu_484_p2;
            lshr_ln702_reg_714 <= lshr_ln702_fu_499_p2;
            or_ln_reg_704[0] <= or_ln_fu_476_p3[0];
            shl_ln702_reg_719 <= shl_ln702_fu_513_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state57)) begin
            lshr_ln702_1_reg_724 <= {{add_ln702_3_fu_534_p2[63:1]}};
            tmp_31_reg_729 <= add_ln702_3_fu_534_p2[32'd54];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state55)) begin
            lshr_ln702_2_reg_699 <= lshr_ln702_2_fu_400_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state53)) begin
            select_ln702_reg_663 <= select_ln702_fu_306_p3;
            tmp_28_reg_658 <= grp_atan2_generic_double_Pipeline_1_fu_128_z_out[32'd85];
            tmp_s_reg_671 <= {{select_ln702_fu_306_p3[85:22]}};
            trunc_ln702_1_reg_677 <= trunc_ln702_1_fu_324_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state54)) begin
            sub_ln702_1_reg_687   <= sub_ln702_1_fu_381_p2;
            trunc_ln702_3_reg_682 <= trunc_ln702_3_fu_377_p1;
            trunc_ln702_4_reg_694 <= trunc_ln702_4_fu_387_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            x_reg_650[84 : 33] <= x_fu_273_p4[84 : 33];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            y_3_reg_645 <= y_3_fu_266_p3;
        end
    end

    assign ap_ST_fsm_state100_blk = 1'b0;

    assign ap_ST_fsm_state101_blk = 1'b0;

    assign ap_ST_fsm_state102_blk = 1'b0;

    assign ap_ST_fsm_state103_blk = 1'b0;

    assign ap_ST_fsm_state104_blk = 1'b0;

    assign ap_ST_fsm_state105_blk = 1'b0;

    assign ap_ST_fsm_state106_blk = 1'b0;

    assign ap_ST_fsm_state107_blk = 1'b0;

    assign ap_ST_fsm_state108_blk = 1'b0;

    assign ap_ST_fsm_state109_blk = 1'b0;

    assign ap_ST_fsm_state10_blk  = 1'b0;

    assign ap_ST_fsm_state110_blk = 1'b0;

    assign ap_ST_fsm_state111_blk = 1'b0;

    assign ap_ST_fsm_state112_blk = 1'b0;

    assign ap_ST_fsm_state113_blk = 1'b0;

    assign ap_ST_fsm_state114_blk = 1'b0;

    assign ap_ST_fsm_state115_blk = 1'b0;

    assign ap_ST_fsm_state116_blk = 1'b0;

    assign ap_ST_fsm_state11_blk  = 1'b0;

    assign ap_ST_fsm_state12_blk  = 1'b0;

    assign ap_ST_fsm_state13_blk  = 1'b0;

    assign ap_ST_fsm_state14_blk  = 1'b0;

    assign ap_ST_fsm_state15_blk  = 1'b0;

    assign ap_ST_fsm_state16_blk  = 1'b0;

    assign ap_ST_fsm_state17_blk  = 1'b0;

    assign ap_ST_fsm_state18_blk  = 1'b0;

    assign ap_ST_fsm_state19_blk  = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    always @(*) begin
        if ((grp_atan2_generic_double_Pipeline_1_fu_128_ap_done == 1'b0)) begin
            ap_ST_fsm_state4_blk = 1'b1;
        end else begin
            ap_ST_fsm_state4_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    assign ap_ST_fsm_state73_blk = 1'b0;

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state75_blk = 1'b0;

    assign ap_ST_fsm_state76_blk = 1'b0;

    assign ap_ST_fsm_state77_blk = 1'b0;

    assign ap_ST_fsm_state78_blk = 1'b0;

    assign ap_ST_fsm_state79_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state80_blk = 1'b0;

    assign ap_ST_fsm_state81_blk = 1'b0;

    assign ap_ST_fsm_state82_blk = 1'b0;

    assign ap_ST_fsm_state83_blk = 1'b0;

    assign ap_ST_fsm_state84_blk = 1'b0;

    assign ap_ST_fsm_state85_blk = 1'b0;

    assign ap_ST_fsm_state86_blk = 1'b0;

    assign ap_ST_fsm_state87_blk = 1'b0;

    assign ap_ST_fsm_state88_blk = 1'b0;

    assign ap_ST_fsm_state89_blk = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state90_blk = 1'b0;

    assign ap_ST_fsm_state91_blk = 1'b0;

    assign ap_ST_fsm_state92_blk = 1'b0;

    assign ap_ST_fsm_state93_blk = 1'b0;

    assign ap_ST_fsm_state94_blk = 1'b0;

    assign ap_ST_fsm_state95_blk = 1'b0;

    assign ap_ST_fsm_state96_blk = 1'b0;

    assign ap_ST_fsm_state97_blk = 1'b0;

    assign ap_ST_fsm_state98_blk = 1'b0;

    assign ap_ST_fsm_state99_blk = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state116) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state116) & (icmp_ln655_reg_618 == 1'd1))) begin
            ap_phi_mux_retval_0_phi_fu_116_p8 = grp_fu_137_p2;
        end else begin
            ap_phi_mux_retval_0_phi_fu_116_p8 = retval_0_reg_112;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state116)) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state116)) begin
            ap_return = ap_phi_mux_retval_0_phi_fu_116_p8;
        end else begin
            ap_return = ap_return_preg;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((icmp_ln662_fu_192_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1) & (icmp_ln655_fu_186_p2 == 1'd0) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state116;
                end else if (((icmp_ln662_fu_192_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1) & (icmp_ln655_fu_186_p2 == 1'd0) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else if (((1'b1 == ap_CS_fsm_state1) & (icmp_ln655_fu_186_p2 == 1'd1) & (ap_start == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_state59;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                if (((grp_atan2_generic_double_Pipeline_1_fu_128_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state4))) begin
                    ap_NS_fsm = ap_ST_fsm_state5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                if (((icmp_ln702_fu_286_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state53))) begin
                    ap_NS_fsm = ap_ST_fsm_state116;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state54;
                end
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state116;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end
            ap_ST_fsm_state78: begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
            ap_ST_fsm_state79: begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end
            ap_ST_fsm_state80: begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
            ap_ST_fsm_state81: begin
                ap_NS_fsm = ap_ST_fsm_state82;
            end
            ap_ST_fsm_state82: begin
                ap_NS_fsm = ap_ST_fsm_state83;
            end
            ap_ST_fsm_state83: begin
                ap_NS_fsm = ap_ST_fsm_state84;
            end
            ap_ST_fsm_state84: begin
                ap_NS_fsm = ap_ST_fsm_state85;
            end
            ap_ST_fsm_state85: begin
                ap_NS_fsm = ap_ST_fsm_state86;
            end
            ap_ST_fsm_state86: begin
                ap_NS_fsm = ap_ST_fsm_state87;
            end
            ap_ST_fsm_state87: begin
                ap_NS_fsm = ap_ST_fsm_state88;
            end
            ap_ST_fsm_state88: begin
                ap_NS_fsm = ap_ST_fsm_state89;
            end
            ap_ST_fsm_state89: begin
                ap_NS_fsm = ap_ST_fsm_state90;
            end
            ap_ST_fsm_state90: begin
                ap_NS_fsm = ap_ST_fsm_state91;
            end
            ap_ST_fsm_state91: begin
                ap_NS_fsm = ap_ST_fsm_state92;
            end
            ap_ST_fsm_state92: begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end
            ap_ST_fsm_state93: begin
                ap_NS_fsm = ap_ST_fsm_state94;
            end
            ap_ST_fsm_state94: begin
                ap_NS_fsm = ap_ST_fsm_state95;
            end
            ap_ST_fsm_state95: begin
                ap_NS_fsm = ap_ST_fsm_state96;
            end
            ap_ST_fsm_state96: begin
                ap_NS_fsm = ap_ST_fsm_state97;
            end
            ap_ST_fsm_state97: begin
                ap_NS_fsm = ap_ST_fsm_state98;
            end
            ap_ST_fsm_state98: begin
                ap_NS_fsm = ap_ST_fsm_state99;
            end
            ap_ST_fsm_state99: begin
                ap_NS_fsm = ap_ST_fsm_state100;
            end
            ap_ST_fsm_state100: begin
                ap_NS_fsm = ap_ST_fsm_state101;
            end
            ap_ST_fsm_state101: begin
                ap_NS_fsm = ap_ST_fsm_state102;
            end
            ap_ST_fsm_state102: begin
                ap_NS_fsm = ap_ST_fsm_state103;
            end
            ap_ST_fsm_state103: begin
                ap_NS_fsm = ap_ST_fsm_state104;
            end
            ap_ST_fsm_state104: begin
                ap_NS_fsm = ap_ST_fsm_state105;
            end
            ap_ST_fsm_state105: begin
                ap_NS_fsm = ap_ST_fsm_state106;
            end
            ap_ST_fsm_state106: begin
                ap_NS_fsm = ap_ST_fsm_state107;
            end
            ap_ST_fsm_state107: begin
                ap_NS_fsm = ap_ST_fsm_state108;
            end
            ap_ST_fsm_state108: begin
                ap_NS_fsm = ap_ST_fsm_state109;
            end
            ap_ST_fsm_state109: begin
                ap_NS_fsm = ap_ST_fsm_state110;
            end
            ap_ST_fsm_state110: begin
                ap_NS_fsm = ap_ST_fsm_state111;
            end
            ap_ST_fsm_state111: begin
                ap_NS_fsm = ap_ST_fsm_state112;
            end
            ap_ST_fsm_state112: begin
                ap_NS_fsm = ap_ST_fsm_state113;
            end
            ap_ST_fsm_state113: begin
                ap_NS_fsm = ap_ST_fsm_state114;
            end
            ap_ST_fsm_state114: begin
                ap_NS_fsm = ap_ST_fsm_state115;
            end
            ap_ST_fsm_state115: begin
                ap_NS_fsm = ap_ST_fsm_state116;
            end
            ap_ST_fsm_state116: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign LD_fu_586_p5 = {{tmp_17_fu_579_p3}, {zext_ln702_3_fu_558_p1[51:0]}};

    assign add_ln655_fu_176_p2 = (zext_ln655_fu_172_p1 + 12'd27);

    assign add_ln702_1_fu_406_p2 = ($signed(sub_ln702_1_reg_687) + $signed(32'd4294967243));

    assign add_ln702_2_fu_490_p2 = ($signed(sub_ln702_1_reg_687) + $signed(32'd4294967242));

    assign add_ln702_3_fu_534_p2 = (select_ln702_2_fu_524_p3 + zext_ln702_2_fu_531_p1);

    assign add_ln702_4_fu_573_p2 = (sub_ln702_3_fu_568_p2 + select_ln702_3_fu_561_p3);

    assign add_ln702_fu_363_p2 = (trunc_ln702_2_fu_359_p1 + trunc_ln702_fu_335_p1);

    assign and_ln702_1_fu_464_p2 = (xor_ln702_fu_451_p2 & bit_select27_i_i_fu_457_p3);

    assign and_ln702_2_fu_427_p2 = (select_ln702_reg_663 & lshr_ln702_2_reg_699);

    assign and_ln702_fu_437_p2 = (icmp_ln702_3_fu_431_p2 & icmp_ln702_2_fu_421_p2);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state116 = ap_CS_fsm[32'd115];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state53 = ap_CS_fsm[32'd52];

    assign ap_CS_fsm_state54 = ap_CS_fsm[32'd53];

    assign ap_CS_fsm_state55 = ap_CS_fsm[32'd54];

    assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];

    assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];

    assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];

    assign bit_select27_i_i_fu_457_p3 = select_ln702_reg_663[add_ln702_1_fu_406_p2];

    assign bitcast_ln753_fu_598_p1 = LD_fu_586_p5;

    assign d_exp_fu_198_p2 = (zext_ln655_1_fu_182_p1 - zext_ln655_fu_172_p1);

    assign data_5_fu_158_p1 = y_in;

    assign data_fu_144_p1 = x_in;

    assign fps_x_exp_fu_148_p4 = {{data_fu_144_p1[62:52]}};

    assign fps_y_exp_fu_162_p4 = {{data_5_fu_158_p1[62:52]}};

    assign grp_atan2_generic_double_Pipeline_1_fu_128_ap_start = grp_atan2_generic_double_Pipeline_1_fu_128_ap_start_reg;

    assign icmp_ln655_fu_186_p2 = ((add_ln655_fu_176_p2 < zext_ln655_1_fu_182_p1) ? 1'b1 : 1'b0);

    assign icmp_ln662_fu_192_p2 = ((fps_y_exp_fu_162_p4 == 11'd0) ? 1'b1 : 1'b0);

    assign icmp_ln702_1_fu_339_p2 = ((tmp_s_reg_671 == 64'd0) ? 1'b1 : 1'b0);

    assign icmp_ln702_2_fu_421_p2 = (($signed(tmp_29_fu_411_p4) > $signed(31'd0)) ? 1'b1 : 1'b0);

    assign icmp_ln702_3_fu_431_p2 = ((and_ln702_2_fu_427_p2 != 86'd0) ? 1'b1 : 1'b0);

    assign icmp_ln702_4_fu_484_p2 = (($signed(
        add_ln702_1_fu_406_p2
    ) > $signed(
        32'd0
    )) ? 1'b1 : 1'b0);

    assign icmp_ln702_fu_286_p2 = ((grp_atan2_generic_double_Pipeline_1_fu_128_z_out == 86'd0) ? 1'b1 : 1'b0);

    assign lshr_ln695_fu_260_p2 = zext_ln681_fu_247_p1 >> zext_ln695_fu_251_p1;

    assign lshr_ln702_2_fu_400_p2 = 86'd77371252455336267181195263 >> zext_ln702_4_fu_396_p1;

    assign lshr_ln702_fu_499_p2 = select_ln702_reg_663 >> zext_ln702_fu_495_p1;

    assign or_ln702_fu_470_p2 = (and_ln702_fu_437_p2 | and_ln702_1_fu_464_p2);

    assign or_ln_fu_476_p3 = {{1'd0}, {or_ln702_fu_470_p2}};

    assign select_ln695_fu_230_p3 = ((tmp_fu_216_p3[0:0] == 1'b1) ? sub_ln695_fu_224_p2 : trunc_ln688_fu_204_p1);

    assign select_ln702_1_fu_369_p3 = ((icmp_ln702_1_fu_339_p2[0:0] == 1'b1) ? add_ln702_fu_363_p2 : trunc_ln702_fu_335_p1);

    assign select_ln702_2_fu_524_p3 = ((icmp_ln702_4_reg_709[0:0] == 1'b1) ? trunc_ln702_5_fu_518_p1 : trunc_ln702_6_fu_521_p1);

    assign select_ln702_3_fu_561_p3 = ((tmp_31_reg_729[0:0] == 1'b1) ? 11'd1023 : 11'd1022);

    assign select_ln702_fu_306_p3 = ((tmp_28_fu_292_p3[0:0] == 1'b1) ? sub_ln702_fu_300_p2 : grp_atan2_generic_double_Pipeline_1_fu_128_z_out);

    assign shl_ln695_fu_254_p2 = zext_ln681_fu_247_p1 << zext_ln695_fu_251_p1;

    assign shl_ln702_fu_513_p2 = select_ln702_reg_663 << zext_ln702_1_fu_509_p1;

    assign sub_ln695_fu_224_p2 = (11'd0 - trunc_ln688_fu_204_p1);

    assign sub_ln702_1_fu_381_p2 = (32'd86 - select_ln702_1_fu_369_p3);

    assign sub_ln702_2_fu_504_p2 = (32'd54 - sub_ln702_1_reg_687);

    assign sub_ln702_3_fu_568_p2 = (11'd1 - trunc_ln702_3_reg_682);

    assign sub_ln702_4_fu_391_p2 = (7'd12 - trunc_ln702_4_reg_694);

    assign sub_ln702_fu_300_p2 = (86'd0 - grp_atan2_generic_double_Pipeline_1_fu_128_z_out);

    always @(tmp_s_reg_671) begin
        if (tmp_s_reg_671[63] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd0;
        end else if (tmp_s_reg_671[62] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd1;
        end else if (tmp_s_reg_671[61] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd2;
        end else if (tmp_s_reg_671[60] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd3;
        end else if (tmp_s_reg_671[59] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd4;
        end else if (tmp_s_reg_671[58] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd5;
        end else if (tmp_s_reg_671[57] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd6;
        end else if (tmp_s_reg_671[56] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd7;
        end else if (tmp_s_reg_671[55] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd8;
        end else if (tmp_s_reg_671[54] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd9;
        end else if (tmp_s_reg_671[53] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd10;
        end else if (tmp_s_reg_671[52] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd11;
        end else if (tmp_s_reg_671[51] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd12;
        end else if (tmp_s_reg_671[50] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd13;
        end else if (tmp_s_reg_671[49] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd14;
        end else if (tmp_s_reg_671[48] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd15;
        end else if (tmp_s_reg_671[47] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd16;
        end else if (tmp_s_reg_671[46] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd17;
        end else if (tmp_s_reg_671[45] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd18;
        end else if (tmp_s_reg_671[44] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd19;
        end else if (tmp_s_reg_671[43] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd20;
        end else if (tmp_s_reg_671[42] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd21;
        end else if (tmp_s_reg_671[41] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd22;
        end else if (tmp_s_reg_671[40] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd23;
        end else if (tmp_s_reg_671[39] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd24;
        end else if (tmp_s_reg_671[38] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd25;
        end else if (tmp_s_reg_671[37] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd26;
        end else if (tmp_s_reg_671[36] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd27;
        end else if (tmp_s_reg_671[35] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd28;
        end else if (tmp_s_reg_671[34] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd29;
        end else if (tmp_s_reg_671[33] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd30;
        end else if (tmp_s_reg_671[32] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd31;
        end else if (tmp_s_reg_671[31] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd32;
        end else if (tmp_s_reg_671[30] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd33;
        end else if (tmp_s_reg_671[29] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd34;
        end else if (tmp_s_reg_671[28] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd35;
        end else if (tmp_s_reg_671[27] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd36;
        end else if (tmp_s_reg_671[26] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd37;
        end else if (tmp_s_reg_671[25] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd38;
        end else if (tmp_s_reg_671[24] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd39;
        end else if (tmp_s_reg_671[23] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd40;
        end else if (tmp_s_reg_671[22] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd41;
        end else if (tmp_s_reg_671[21] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd42;
        end else if (tmp_s_reg_671[20] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd43;
        end else if (tmp_s_reg_671[19] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd44;
        end else if (tmp_s_reg_671[18] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd45;
        end else if (tmp_s_reg_671[17] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd46;
        end else if (tmp_s_reg_671[16] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd47;
        end else if (tmp_s_reg_671[15] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd48;
        end else if (tmp_s_reg_671[14] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd49;
        end else if (tmp_s_reg_671[13] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd50;
        end else if (tmp_s_reg_671[12] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd51;
        end else if (tmp_s_reg_671[11] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd52;
        end else if (tmp_s_reg_671[10] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd53;
        end else if (tmp_s_reg_671[9] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd54;
        end else if (tmp_s_reg_671[8] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd55;
        end else if (tmp_s_reg_671[7] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd56;
        end else if (tmp_s_reg_671[6] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd57;
        end else if (tmp_s_reg_671[5] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd58;
        end else if (tmp_s_reg_671[4] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd59;
        end else if (tmp_s_reg_671[3] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd60;
        end else if (tmp_s_reg_671[2] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd61;
        end else if (tmp_s_reg_671[1] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd62;
        end else if (tmp_s_reg_671[0] == 1'b1) begin
            tmp_12_fu_328_p3 = 64'd63;
        end else begin
            tmp_12_fu_328_p3 = 64'd64;
        end
    end

    assign tmp_14_fu_344_p3 = {{trunc_ln702_1_reg_677}, {42'd4398046511103}};

    always @(tmp_14_fu_344_p3) begin
        if (tmp_14_fu_344_p3[63] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd0;
        end else if (tmp_14_fu_344_p3[62] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd1;
        end else if (tmp_14_fu_344_p3[61] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd2;
        end else if (tmp_14_fu_344_p3[60] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd3;
        end else if (tmp_14_fu_344_p3[59] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd4;
        end else if (tmp_14_fu_344_p3[58] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd5;
        end else if (tmp_14_fu_344_p3[57] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd6;
        end else if (tmp_14_fu_344_p3[56] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd7;
        end else if (tmp_14_fu_344_p3[55] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd8;
        end else if (tmp_14_fu_344_p3[54] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd9;
        end else if (tmp_14_fu_344_p3[53] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd10;
        end else if (tmp_14_fu_344_p3[52] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd11;
        end else if (tmp_14_fu_344_p3[51] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd12;
        end else if (tmp_14_fu_344_p3[50] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd13;
        end else if (tmp_14_fu_344_p3[49] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd14;
        end else if (tmp_14_fu_344_p3[48] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd15;
        end else if (tmp_14_fu_344_p3[47] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd16;
        end else if (tmp_14_fu_344_p3[46] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd17;
        end else if (tmp_14_fu_344_p3[45] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd18;
        end else if (tmp_14_fu_344_p3[44] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd19;
        end else if (tmp_14_fu_344_p3[43] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd20;
        end else if (tmp_14_fu_344_p3[42] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd21;
        end else if (tmp_14_fu_344_p3[41] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd22;
        end else if (tmp_14_fu_344_p3[40] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd23;
        end else if (tmp_14_fu_344_p3[39] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd24;
        end else if (tmp_14_fu_344_p3[38] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd25;
        end else if (tmp_14_fu_344_p3[37] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd26;
        end else if (tmp_14_fu_344_p3[36] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd27;
        end else if (tmp_14_fu_344_p3[35] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd28;
        end else if (tmp_14_fu_344_p3[34] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd29;
        end else if (tmp_14_fu_344_p3[33] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd30;
        end else if (tmp_14_fu_344_p3[32] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd31;
        end else if (tmp_14_fu_344_p3[31] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd32;
        end else if (tmp_14_fu_344_p3[30] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd33;
        end else if (tmp_14_fu_344_p3[29] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd34;
        end else if (tmp_14_fu_344_p3[28] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd35;
        end else if (tmp_14_fu_344_p3[27] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd36;
        end else if (tmp_14_fu_344_p3[26] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd37;
        end else if (tmp_14_fu_344_p3[25] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd38;
        end else if (tmp_14_fu_344_p3[24] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd39;
        end else if (tmp_14_fu_344_p3[23] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd40;
        end else if (tmp_14_fu_344_p3[22] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd41;
        end else if (tmp_14_fu_344_p3[21] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd42;
        end else if (tmp_14_fu_344_p3[20] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd43;
        end else if (tmp_14_fu_344_p3[19] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd44;
        end else if (tmp_14_fu_344_p3[18] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd45;
        end else if (tmp_14_fu_344_p3[17] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd46;
        end else if (tmp_14_fu_344_p3[16] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd47;
        end else if (tmp_14_fu_344_p3[15] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd48;
        end else if (tmp_14_fu_344_p3[14] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd49;
        end else if (tmp_14_fu_344_p3[13] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd50;
        end else if (tmp_14_fu_344_p3[12] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd51;
        end else if (tmp_14_fu_344_p3[11] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd52;
        end else if (tmp_14_fu_344_p3[10] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd53;
        end else if (tmp_14_fu_344_p3[9] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd54;
        end else if (tmp_14_fu_344_p3[8] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd55;
        end else if (tmp_14_fu_344_p3[7] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd56;
        end else if (tmp_14_fu_344_p3[6] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd57;
        end else if (tmp_14_fu_344_p3[5] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd58;
        end else if (tmp_14_fu_344_p3[4] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd59;
        end else if (tmp_14_fu_344_p3[3] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd60;
        end else if (tmp_14_fu_344_p3[2] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd61;
        end else if (tmp_14_fu_344_p3[1] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd62;
        end else if (tmp_14_fu_344_p3[0] == 1'b1) begin
            tmp_15_fu_351_p3 = 64'd63;
        end else begin
            tmp_15_fu_351_p3 = 64'd64;
        end
    end

    assign tmp_17_fu_579_p3 = {{tmp_28_reg_658}, {add_ln702_4_fu_573_p2}};

    assign tmp_28_fu_292_p3 = grp_atan2_generic_double_Pipeline_1_fu_128_z_out[32'd85];

    assign tmp_29_fu_411_p4 = {{add_ln702_1_fu_406_p2[31:1]}};

    assign tmp_30_fu_443_p3 = add_ln702_1_fu_406_p2[32'd31];

    assign tmp_fu_216_p3 = d_exp_fu_198_p2[32'd11];

    assign trunc_ln505_2_fu_212_p1 = data_5_fu_158_p1[51:0];

    assign trunc_ln505_fu_208_p1 = data_fu_144_p1[51:0];

    assign trunc_ln688_fu_204_p1 = d_exp_fu_198_p2[10:0];

    assign trunc_ln702_1_fu_324_p1 = select_ln702_fu_306_p3[21:0];

    assign trunc_ln702_2_fu_359_p1 = tmp_15_fu_351_p3[31:0];

    assign trunc_ln702_3_fu_377_p1 = select_ln702_1_fu_369_p3[10:0];

    assign trunc_ln702_4_fu_387_p1 = sub_ln702_1_fu_381_p2[6:0];

    assign trunc_ln702_5_fu_518_p1 = lshr_ln702_reg_714[63:0];

    assign trunc_ln702_6_fu_521_p1 = shl_ln702_reg_719[63:0];

    assign trunc_ln702_fu_335_p1 = tmp_12_fu_328_p3[31:0];

    assign x_fu_273_p4 = {{{{1'd1}, {trunc_ln505_reg_625}}}, {33'd0}};

    assign xor_ln702_fu_451_p2 = (tmp_30_fu_443_p3 ^ 1'd1);

    assign y_3_fu_266_p3 = ((tmp_reg_635[0:0] == 1'b1) ? shl_ln695_fu_254_p2 : lshr_ln695_fu_260_p2);

    assign y_fu_238_p4 = {{{{1'd1}, {trunc_ln505_2_reg_630}}}, {33'd0}};

    assign zext_ln655_1_fu_182_p1 = fps_x_exp_fu_148_p4;

    assign zext_ln655_fu_172_p1 = fps_y_exp_fu_162_p4;

    assign zext_ln681_fu_247_p1 = y_fu_238_p4;

    assign zext_ln695_fu_251_p1 = select_ln695_reg_640;

    assign zext_ln702_1_fu_509_p1 = sub_ln702_2_fu_504_p2;

    assign zext_ln702_2_fu_531_p1 = or_ln_reg_704;

    assign zext_ln702_3_fu_558_p1 = lshr_ln702_1_reg_724;

    assign zext_ln702_4_fu_396_p1 = sub_ln702_4_fu_391_p2;

    assign zext_ln702_fu_495_p1 = add_ln702_2_fu_490_p2;

    always @(posedge ap_clk) begin
        x_reg_650[32:0] <= 33'b000000000000000000000000000000000;
        x_reg_650[85] <= 1'b1;
        or_ln_reg_704[1] <= 1'b0;
    end

endmodule  //main_atan2_generic_double_s
