/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns / 1ps

module main_dcmp_64ns_64ns_1_2_no_dsp_1_x #(
    parameter ID         = 1,
              NUM_STAGE  = 2,
              din0_WIDTH = 32,
              din1_WIDTH = 32,
              dout_WIDTH = 1
) (
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  ce,
    input  wire [din0_WIDTH-1:0] din0,
    input  wire [din1_WIDTH-1:0] din1,
    input  wire [           4:0] opcode,
    output wire [dout_WIDTH-1:0] dout
);
    //------------------------Parameter----------------------
    // AutoESL opcode
    localparam [4:0]
    AP_OEQ = 5'b00001,
    AP_OGT = 5'b00010,
    AP_OGE = 5'b00011,
    AP_OLT = 5'b00100,
    AP_OLE = 5'b00101,
    AP_ONE = 5'b00110,
    AP_UNO = 5'b01000;
    // FPV6 opcode
    localparam [7:0]
    OP_EQ = 8'b00010100,
    OP_GT = 8'b00100100,
    OP_GE = 8'b00110100,
    OP_LT = 8'b00001100,
    OP_LE = 8'b00011100,
    OP_NE = 8'b00101100,
    OP_UO = 8'b00000100;
    //------------------------Local signal-------------------
    wire                  a_tvalid;
    wire [din0_WIDTH-1:0] a_tdata;
    wire                  b_tvalid;
    wire [din1_WIDTH-1:0] b_tdata;
    wire                  op_tvalid;
    reg  [           7:0] op_tdata;
    wire                  r_tvalid;
    wire [           7:0] r_tdata;
    reg  [din0_WIDTH-1:0] din0_buf1;
    reg  [din1_WIDTH-1:0] din1_buf1;
    reg  [           4:0] opcode_buf1;
    reg                   ce_r;
    wire [dout_WIDTH-1:0] dout_i;
    reg  [dout_WIDTH-1:0] dout_r;
    //------------------------Instantiation------------------
    main_dcmp_64ns_64ns_1_2_no_dsp_1_x_ip main_dcmp_64ns_64ns_1_2_no_dsp_1_x_ip_u (
        .s_axis_a_tvalid        (a_tvalid),
        .s_axis_a_tdata         (a_tdata),
        .s_axis_b_tvalid        (b_tvalid),
        .s_axis_b_tdata         (b_tdata),
        .s_axis_operation_tvalid(op_tvalid),
        .s_axis_operation_tdata (op_tdata),
        .m_axis_result_tvalid   (r_tvalid),
        .m_axis_result_tdata    (r_tdata)
    );
    //------------------------Body---------------------------
    assign a_tvalid  = 1'b1;
    assign a_tdata   = din0_buf1;
    assign b_tvalid  = 1'b1;
    assign b_tdata   = din1_buf1;
    assign op_tvalid = 1'b1;
    assign dout_i    = r_tdata[0];

    always @(*) begin
        case (opcode_buf1)
            AP_OEQ:  op_tdata = OP_EQ;
            AP_OGT:  op_tdata = OP_GT;
            AP_OGE:  op_tdata = OP_GE;
            AP_OLT:  op_tdata = OP_LT;
            AP_OLE:  op_tdata = OP_LE;
            AP_ONE:  op_tdata = OP_NE;
            AP_UNO:  op_tdata = OP_UO;
            default: op_tdata = OP_EQ;
        endcase
    end

    always @(posedge clk) begin
        if (ce) begin
            din0_buf1   <= din0;
            din1_buf1   <= din1;
            opcode_buf1 <= opcode;
        end
    end

    always @(posedge clk) begin
        ce_r <= ce;
    end

    always @(posedge clk) begin
        if (ce_r) begin
            dout_r <= dout_i;
        end
    end

    assign dout = ce_r ? dout_i : dout_r;
endmodule
