/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_rayCast_Pipeline_VITIS_LOOP_222_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    xRay,
    yRay,
    step,
    xStep,
    yStep,
    tmp_30,
    trunc_ln230_1,
    empty,
    pf_address0,
    pf_ce0,
    pf_q0,
    pf_load_6,
    trunc_ln235_3,
    bitcast_ln235,
    dist_1_out,
    dist_1_out_ap_vld,
    grp_fu_427_p_din0,
    grp_fu_427_p_dout0,
    grp_fu_427_p_ce,
    grp_fu_430_p_din0,
    grp_fu_430_p_din1,
    grp_fu_430_p_opcode,
    grp_fu_430_p_dout0,
    grp_fu_430_p_ce,
    grp_fu_179_p_din0,
    grp_fu_179_p_din1,
    grp_fu_179_p_opcode,
    grp_fu_179_p_dout0,
    grp_fu_179_p_ce,
    grp_fu_434_p_din0,
    grp_fu_434_p_din1,
    grp_fu_434_p_dout0,
    grp_fu_434_p_ce,
    grp_fu_438_p_din0,
    grp_fu_438_p_din1,
    grp_fu_438_p_opcode,
    grp_fu_438_p_dout0,
    grp_fu_438_p_ce
);

    parameter ap_ST_fsm_state1 = 82'd1;
    parameter ap_ST_fsm_state2 = 82'd2;
    parameter ap_ST_fsm_state3 = 82'd4;
    parameter ap_ST_fsm_state4 = 82'd8;
    parameter ap_ST_fsm_state5 = 82'd16;
    parameter ap_ST_fsm_state6 = 82'd32;
    parameter ap_ST_fsm_state7 = 82'd64;
    parameter ap_ST_fsm_state8 = 82'd128;
    parameter ap_ST_fsm_state9 = 82'd256;
    parameter ap_ST_fsm_state10 = 82'd512;
    parameter ap_ST_fsm_state11 = 82'd1024;
    parameter ap_ST_fsm_state12 = 82'd2048;
    parameter ap_ST_fsm_state13 = 82'd4096;
    parameter ap_ST_fsm_state14 = 82'd8192;
    parameter ap_ST_fsm_state15 = 82'd16384;
    parameter ap_ST_fsm_state16 = 82'd32768;
    parameter ap_ST_fsm_state17 = 82'd65536;
    parameter ap_ST_fsm_state18 = 82'd131072;
    parameter ap_ST_fsm_state19 = 82'd262144;
    parameter ap_ST_fsm_state20 = 82'd524288;
    parameter ap_ST_fsm_state21 = 82'd1048576;
    parameter ap_ST_fsm_state22 = 82'd2097152;
    parameter ap_ST_fsm_state23 = 82'd4194304;
    parameter ap_ST_fsm_state24 = 82'd8388608;
    parameter ap_ST_fsm_state25 = 82'd16777216;
    parameter ap_ST_fsm_state26 = 82'd33554432;
    parameter ap_ST_fsm_state27 = 82'd67108864;
    parameter ap_ST_fsm_state28 = 82'd134217728;
    parameter ap_ST_fsm_state29 = 82'd268435456;
    parameter ap_ST_fsm_state30 = 82'd536870912;
    parameter ap_ST_fsm_state31 = 82'd1073741824;
    parameter ap_ST_fsm_state32 = 82'd2147483648;
    parameter ap_ST_fsm_state33 = 82'd4294967296;
    parameter ap_ST_fsm_state34 = 82'd8589934592;
    parameter ap_ST_fsm_state35 = 82'd17179869184;
    parameter ap_ST_fsm_state36 = 82'd34359738368;
    parameter ap_ST_fsm_state37 = 82'd68719476736;
    parameter ap_ST_fsm_state38 = 82'd137438953472;
    parameter ap_ST_fsm_state39 = 82'd274877906944;
    parameter ap_ST_fsm_state40 = 82'd549755813888;
    parameter ap_ST_fsm_state41 = 82'd1099511627776;
    parameter ap_ST_fsm_state42 = 82'd2199023255552;
    parameter ap_ST_fsm_state43 = 82'd4398046511104;
    parameter ap_ST_fsm_state44 = 82'd8796093022208;
    parameter ap_ST_fsm_state45 = 82'd17592186044416;
    parameter ap_ST_fsm_state46 = 82'd35184372088832;
    parameter ap_ST_fsm_state47 = 82'd70368744177664;
    parameter ap_ST_fsm_state48 = 82'd140737488355328;
    parameter ap_ST_fsm_state49 = 82'd281474976710656;
    parameter ap_ST_fsm_state50 = 82'd562949953421312;
    parameter ap_ST_fsm_state51 = 82'd1125899906842624;
    parameter ap_ST_fsm_state52 = 82'd2251799813685248;
    parameter ap_ST_fsm_state53 = 82'd4503599627370496;
    parameter ap_ST_fsm_state54 = 82'd9007199254740992;
    parameter ap_ST_fsm_state55 = 82'd18014398509481984;
    parameter ap_ST_fsm_state56 = 82'd36028797018963968;
    parameter ap_ST_fsm_state57 = 82'd72057594037927936;
    parameter ap_ST_fsm_state58 = 82'd144115188075855872;
    parameter ap_ST_fsm_state59 = 82'd288230376151711744;
    parameter ap_ST_fsm_state60 = 82'd576460752303423488;
    parameter ap_ST_fsm_state61 = 82'd1152921504606846976;
    parameter ap_ST_fsm_state62 = 82'd2305843009213693952;
    parameter ap_ST_fsm_state63 = 82'd4611686018427387904;
    parameter ap_ST_fsm_state64 = 82'd9223372036854775808;
    parameter ap_ST_fsm_state65 = 82'd18446744073709551616;
    parameter ap_ST_fsm_state66 = 82'd36893488147419103232;
    parameter ap_ST_fsm_state67 = 82'd73786976294838206464;
    parameter ap_ST_fsm_state68 = 82'd147573952589676412928;
    parameter ap_ST_fsm_state69 = 82'd295147905179352825856;
    parameter ap_ST_fsm_state70 = 82'd590295810358705651712;
    parameter ap_ST_fsm_state71 = 82'd1180591620717411303424;
    parameter ap_ST_fsm_state72 = 82'd2361183241434822606848;
    parameter ap_ST_fsm_state73 = 82'd4722366482869645213696;
    parameter ap_ST_fsm_state74 = 82'd9444732965739290427392;
    parameter ap_ST_fsm_state75 = 82'd18889465931478580854784;
    parameter ap_ST_fsm_state76 = 82'd37778931862957161709568;
    parameter ap_ST_fsm_state77 = 82'd75557863725914323419136;
    parameter ap_ST_fsm_state78 = 82'd151115727451828646838272;
    parameter ap_ST_fsm_state79 = 82'd302231454903657293676544;
    parameter ap_ST_fsm_state80 = 82'd604462909807314587353088;
    parameter ap_ST_fsm_state81 = 82'd1208925819614629174706176;
    parameter ap_ST_fsm_state82 = 82'd2417851639229258349412352;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] xRay;
    input [63:0] yRay;
    input [63:0] step;
    input [63:0] xStep;
    input [63:0] yStep;
    input [10:0] tmp_30;
    input [51:0] trunc_ln230_1;
    input [63:0] empty;
    output [16:0] pf_address0;
    output pf_ce0;
    input [255:0] pf_q0;
    input [190:0] pf_load_6;
    input [51:0] trunc_ln235_3;
    input [63:0] bitcast_ln235;
    output [63:0] dist_1_out;
    output dist_1_out_ap_vld;
    output [31:0] grp_fu_427_p_din0;
    input [63:0] grp_fu_427_p_dout0;
    output grp_fu_427_p_ce;
    output [31:0] grp_fu_430_p_din0;
    output [31:0] grp_fu_430_p_din1;
    output [4:0] grp_fu_430_p_opcode;
    input [0:0] grp_fu_430_p_dout0;
    output grp_fu_430_p_ce;
    output [63:0] grp_fu_179_p_din0;
    output [63:0] grp_fu_179_p_din1;
    output [0:0] grp_fu_179_p_opcode;
    input [63:0] grp_fu_179_p_dout0;
    output grp_fu_179_p_ce;
    output [63:0] grp_fu_434_p_din0;
    output [63:0] grp_fu_434_p_din1;
    input [63:0] grp_fu_434_p_dout0;
    output grp_fu_434_p_ce;
    output [63:0] grp_fu_438_p_din0;
    output [63:0] grp_fu_438_p_din1;
    output [4:0] grp_fu_438_p_opcode;
    input [0:0] grp_fu_438_p_dout0;
    output grp_fu_438_p_ce;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg pf_ce0;
    reg dist_1_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [81:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    wire    ap_CS_fsm_state2;
    wire   [0:0] icmp_ln230_4_fu_269_p2;
    reg   [0:0] icmp_ln230_4_reg_916;
    wire   [0:0] icmp_ln230_5_fu_274_p2;
    reg   [0:0] icmp_ln230_5_reg_921;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    reg   [63:0] yRay_2_reg_936;
    wire    ap_CS_fsm_state8;
    reg   [63:0] xRay_2_reg_942;
    wire    ap_CS_fsm_state9;
    reg   [63:0] dist_1_reg_948;
    wire    ap_CS_fsm_state10;
    reg   [0:0] tmp_25_reg_956;
    wire    ap_CS_fsm_state12;
    reg   [0:0] xs_sign_1_reg_961;
    wire    ap_CS_fsm_state67;
    wire   [51:0] trunc_ln505_1_fu_309_p1;
    reg   [51:0] trunc_ln505_1_reg_966;
    wire   [0:0] tmp_24_fu_323_p3;
    reg   [0:0] tmp_24_reg_971;
    wire   [11:0] select_ln18_2_fu_341_p3;
    reg   [11:0] select_ln18_2_reg_976;
    reg   [0:0] xs_sign_reg_981;
    wire    ap_CS_fsm_state68;
    wire   [51:0] trunc_ln505_fu_371_p1;
    reg   [51:0] trunc_ln505_reg_986;
    wire   [0:0] tmp_22_fu_385_p3;
    reg   [0:0] tmp_22_reg_991;
    wire   [11:0] select_ln18_fu_403_p3;
    reg   [11:0] select_ln18_reg_996;
    wire   [31:0] val_1_fu_463_p3;
    reg   [31:0] val_1_reg_1001;
    wire   [31:0] val_fu_522_p3;
    reg   [31:0] val_reg_1007;
    wire    ap_CS_fsm_state69;
    wire   [31:0] result_4_fu_529_p2;
    reg   [31:0] result_4_reg_1013;
    wire   [0:0] or_ln230_2_fu_632_p2;
    reg   [0:0] or_ln230_2_reg_1018;
    wire    ap_CS_fsm_state70;
    wire   [9:0] trunc_ln234_1_fu_646_p1;
    reg   [9:0] trunc_ln234_1_reg_1027;
    wire   [0:0] icmp_ln235_4_fu_659_p2;
    reg   [0:0] icmp_ln235_4_reg_1032;
    wire   [0:0] icmp_ln235_5_fu_665_p2;
    reg   [0:0] icmp_ln235_5_reg_1037;
    wire    ap_CS_fsm_state72;
    wire    ap_CS_fsm_state73;
    wire   [4:0] trunc_ln234_2_fu_705_p1;
    reg   [4:0] trunc_ln234_2_reg_1052;
    reg   [255:0] pf_load_reg_1057;
    wire    ap_CS_fsm_state74;
    wire   [31:0] trunc_ln234_3_fu_724_p1;
    reg   [31:0] trunc_ln234_3_reg_1062;
    wire    ap_CS_fsm_state75;
    wire   [0:0] icmp_ln235_fu_742_p2;
    reg   [0:0] icmp_ln235_reg_1067;
    wire   [0:0] icmp_ln235_1_fu_748_p2;
    reg   [0:0] icmp_ln235_1_reg_1072;
    wire   [31:0] bitcast_ln234_fu_754_p1;
    reg   [63:0] occ_reg_1083;
    wire    ap_CS_fsm_state77;
    reg   [0:0] tmp_28_reg_1089;
    wire   [0:0] icmp_ln235_2_fu_776_p2;
    reg   [0:0] icmp_ln235_2_reg_1094;
    wire    ap_CS_fsm_state78;
    wire   [0:0] icmp_ln235_3_fu_782_p2;
    reg   [0:0] icmp_ln235_3_reg_1099;
    wire   [0:0] and_ln235_2_fu_802_p2;
    reg   [0:0] and_ln235_2_reg_1104;
    wire    ap_CS_fsm_state79;
    wire   [63:0] zext_ln234_3_fu_700_p1;
    reg   [63:0] dist_fu_132;
    wire    ap_CS_fsm_state80;
    wire   [0:0] or_ln235_3_fu_817_p2;
    reg   [63:0] yRay_1_fu_136;
    reg   [63:0] xRay_1_fu_140;
    wire    ap_CS_fsm_state81;
    wire    ap_CS_fsm_state82;
    reg   [63:0] grp_fu_238_p0;
    reg   [63:0] grp_fu_238_p1;
    reg   [63:0] grp_fu_242_p0;
    reg   [63:0] grp_fu_246_p0;
    reg   [63:0] grp_fu_246_p1;
    wire    ap_CS_fsm_state11;
    wire   [63:0] data_4_fu_287_p1;
    wire   [10:0] xs_exp_1_fu_299_p4;
    wire   [11:0] zext_ln486_1_fu_313_p1;
    wire   [11:0] add_ln486_1_fu_317_p2;
    wire   [10:0] sub_ln18_1_fu_331_p2;
    wire  signed [11:0] sext_ln18_2_fu_337_p1;
    wire   [63:0] data_fu_349_p1;
    wire   [10:0] xs_exp_fu_361_p4;
    wire   [11:0] zext_ln486_fu_375_p1;
    wire   [11:0] add_ln486_fu_379_p2;
    wire   [10:0] sub_ln18_fu_393_p2;
    wire  signed [11:0] sext_ln18_fu_399_p1;
    wire   [53:0] mantissa_1_fu_411_p4;
    wire  signed [31:0] sext_ln18_3_fu_424_p1;
    wire   [136:0] zext_ln15_1_fu_420_p1;
    wire   [136:0] zext_ln18_1_fu_427_p1;
    wire   [136:0] lshr_ln18_1_fu_431_p2;
    wire   [136:0] shl_ln18_1_fu_437_p2;
    wire   [31:0] tmp_16_fu_443_p4;
    wire   [31:0] tmp_17_fu_453_p4;
    wire   [53:0] mantissa_fu_470_p4;
    wire  signed [31:0] sext_ln18_1_fu_483_p1;
    wire   [136:0] zext_ln15_fu_479_p1;
    wire   [136:0] zext_ln18_fu_486_p1;
    wire   [136:0] lshr_ln18_fu_490_p2;
    wire   [136:0] shl_ln18_fu_496_p2;
    wire   [31:0] tmp_14_fu_502_p4;
    wire   [31:0] tmp_15_fu_512_p4;
    wire   [31:0] result_1_fu_534_p2;
    wire   [63:0] bitcast_ln230_fu_550_p1;
    wire   [10:0] tmp_s_fu_553_p4;
    wire   [51:0] trunc_ln230_fu_563_p1;
    wire   [0:0] icmp_ln230_3_fu_573_p2;
    wire   [0:0] icmp_ln230_1_fu_567_p2;
    wire   [0:0] or_ln230_fu_579_p2;
    wire   [0:0] or_ln230_1_fu_585_p2;
    wire   [0:0] and_ln230_fu_589_p2;
    wire   [31:0] result_6_fu_545_p3;
    wire   [31:0] result_fu_539_p3;
    wire   [0:0] and_ln230_1_fu_595_p2;
    wire   [0:0] icmp_ln230_fu_600_p2;
    wire   [0:0] icmp_ln230_2_fu_614_p2;
    wire   [0:0] tmp_26_fu_606_p3;
    wire   [0:0] or_ln230_3_fu_626_p2;
    wire   [0:0] or_ln230_4_fu_620_p2;
    wire   [9:0] trunc_ln234_fu_638_p1;
    wire   [10:0] tmp_31_fu_650_p4;
    wire   [11:0] shl_ln_fu_670_p3;
    wire   [14:0] zext_ln234_1_fu_677_p1;
    wire   [14:0] add_ln234_fu_681_p2;
    wire   [21:0] grp_fu_834_p3;
    wire   [16:0] lshr_ln234_1_fu_691_p4;
    wire   [7:0] shl_ln234_1_fu_708_p3;
    wire   [255:0] zext_ln234_4_fu_715_p1;
    wire   [255:0] lshr_ln234_fu_719_p2;
    wire   [7:0] tmp_27_fu_728_p4;
    wire   [22:0] trunc_ln235_fu_738_p1;
    wire   [63:0] bitcast_ln235_1_fu_759_p1;
    wire   [10:0] tmp_29_fu_762_p4;
    wire   [51:0] trunc_ln235_1_fu_772_p1;
    wire   [0:0] or_ln235_1_fu_788_p2;
    wire   [0:0] or_ln235_2_fu_792_p2;
    wire   [0:0] and_ln235_1_fu_796_p2;
    wire   [0:0] or_ln235_fu_808_p2;
    wire   [0:0] and_ln235_fu_812_p2;
    wire   [9:0] grp_fu_834_p0;
    wire   [11:0] grp_fu_834_p1;
    wire   [14:0] grp_fu_834_p2;
    reg   [81:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    wire    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    wire    ap_ST_fsm_state4_blk;
    wire    ap_ST_fsm_state5_blk;
    wire    ap_ST_fsm_state6_blk;
    wire    ap_ST_fsm_state7_blk;
    wire    ap_ST_fsm_state8_blk;
    wire    ap_ST_fsm_state9_blk;
    wire    ap_ST_fsm_state10_blk;
    wire    ap_ST_fsm_state11_blk;
    wire    ap_ST_fsm_state12_blk;
    wire    ap_ST_fsm_state13_blk;
    wire    ap_ST_fsm_state14_blk;
    wire    ap_ST_fsm_state15_blk;
    wire    ap_ST_fsm_state16_blk;
    wire    ap_ST_fsm_state17_blk;
    wire    ap_ST_fsm_state18_blk;
    wire    ap_ST_fsm_state19_blk;
    wire    ap_ST_fsm_state20_blk;
    wire    ap_ST_fsm_state21_blk;
    wire    ap_ST_fsm_state22_blk;
    wire    ap_ST_fsm_state23_blk;
    wire    ap_ST_fsm_state24_blk;
    wire    ap_ST_fsm_state25_blk;
    wire    ap_ST_fsm_state26_blk;
    wire    ap_ST_fsm_state27_blk;
    wire    ap_ST_fsm_state28_blk;
    wire    ap_ST_fsm_state29_blk;
    wire    ap_ST_fsm_state30_blk;
    wire    ap_ST_fsm_state31_blk;
    wire    ap_ST_fsm_state32_blk;
    wire    ap_ST_fsm_state33_blk;
    wire    ap_ST_fsm_state34_blk;
    wire    ap_ST_fsm_state35_blk;
    wire    ap_ST_fsm_state36_blk;
    wire    ap_ST_fsm_state37_blk;
    wire    ap_ST_fsm_state38_blk;
    wire    ap_ST_fsm_state39_blk;
    wire    ap_ST_fsm_state40_blk;
    wire    ap_ST_fsm_state41_blk;
    wire    ap_ST_fsm_state42_blk;
    wire    ap_ST_fsm_state43_blk;
    wire    ap_ST_fsm_state44_blk;
    wire    ap_ST_fsm_state45_blk;
    wire    ap_ST_fsm_state46_blk;
    wire    ap_ST_fsm_state47_blk;
    wire    ap_ST_fsm_state48_blk;
    wire    ap_ST_fsm_state49_blk;
    wire    ap_ST_fsm_state50_blk;
    wire    ap_ST_fsm_state51_blk;
    wire    ap_ST_fsm_state52_blk;
    wire    ap_ST_fsm_state53_blk;
    wire    ap_ST_fsm_state54_blk;
    wire    ap_ST_fsm_state55_blk;
    wire    ap_ST_fsm_state56_blk;
    wire    ap_ST_fsm_state57_blk;
    wire    ap_ST_fsm_state58_blk;
    wire    ap_ST_fsm_state59_blk;
    wire    ap_ST_fsm_state60_blk;
    wire    ap_ST_fsm_state61_blk;
    wire    ap_ST_fsm_state62_blk;
    wire    ap_ST_fsm_state63_blk;
    wire    ap_ST_fsm_state64_blk;
    wire    ap_ST_fsm_state65_blk;
    wire    ap_ST_fsm_state66_blk;
    wire    ap_ST_fsm_state67_blk;
    wire    ap_ST_fsm_state68_blk;
    wire    ap_ST_fsm_state69_blk;
    wire    ap_ST_fsm_state70_blk;
    wire    ap_ST_fsm_state71_blk;
    wire    ap_ST_fsm_state72_blk;
    wire    ap_ST_fsm_state73_blk;
    wire    ap_ST_fsm_state74_blk;
    wire    ap_ST_fsm_state75_blk;
    wire    ap_ST_fsm_state76_blk;
    wire    ap_ST_fsm_state77_blk;
    wire    ap_ST_fsm_state78_blk;
    wire    ap_ST_fsm_state79_blk;
    wire    ap_ST_fsm_state80_blk;
    wire    ap_ST_fsm_state81_blk;
    wire    ap_ST_fsm_state82_blk;
    wire   [21:0] grp_fu_834_p00;
    wire   [21:0] grp_fu_834_p20;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 82'd1;
        #0 dist_fu_132 = 64'd0;
        #0 yRay_1_fu_136 = 64'd0;
        #0 xRay_1_fu_140 = 64'd0;
    end

    main_mac_muladd_10ns_12ns_15ns_22_4_1 #(
        .ID(1),
        .NUM_STAGE(4),
        .din0_WIDTH(10),
        .din1_WIDTH(12),
        .din2_WIDTH(15),
        .dout_WIDTH(22)
    ) mac_muladd_10ns_12ns_15ns_22_4_1_U142 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_834_p0),
        .din1(grp_fu_834_p1),
        .din2(grp_fu_834_p2),
        .ce(1'b1),
        .dout(grp_fu_834_p3)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            dist_fu_132 <= 64'd0;
        end else if (((or_ln235_3_fu_817_p2 == 1'd0) & (or_ln230_2_reg_1018 == 1'd0) & (1'b1 == ap_CS_fsm_state80))) begin
            dist_fu_132 <= dist_1_reg_948;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            xRay_1_fu_140 <= xRay;
        end else if (((or_ln235_3_fu_817_p2 == 1'd0) & (or_ln230_2_reg_1018 == 1'd0) & (1'b1 == ap_CS_fsm_state80))) begin
            xRay_1_fu_140 <= xRay_2_reg_942;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            yRay_1_fu_136 <= yRay;
        end else if (((or_ln235_3_fu_817_p2 == 1'd0) & (or_ln230_2_reg_1018 == 1'd0) & (1'b1 == ap_CS_fsm_state80))) begin
            yRay_1_fu_136 <= yRay_2_reg_936;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state79)) begin
            and_ln235_2_reg_1104 <= and_ln235_2_fu_802_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            dist_1_reg_948 <= grp_fu_179_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            icmp_ln230_4_reg_916 <= icmp_ln230_4_fu_269_p2;
            icmp_ln230_5_reg_921 <= icmp_ln230_5_fu_274_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state75)) begin
            icmp_ln235_1_reg_1072 <= icmp_ln235_1_fu_748_p2;
            icmp_ln235_reg_1067 <= icmp_ln235_fu_742_p2;
            trunc_ln234_3_reg_1062 <= trunc_ln234_3_fu_724_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state78)) begin
            icmp_ln235_2_reg_1094 <= icmp_ln235_2_fu_776_p2;
            icmp_ln235_3_reg_1099 <= icmp_ln235_3_fu_782_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state70)) begin
            icmp_ln235_4_reg_1032 <= icmp_ln235_4_fu_659_p2;
            icmp_ln235_5_reg_1037 <= icmp_ln235_5_fu_665_p2;
            or_ln230_2_reg_1018 <= or_ln230_2_fu_632_p2;
            trunc_ln234_1_reg_1027 <= trunc_ln234_1_fu_646_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state77)) begin
            occ_reg_1083 <= grp_fu_427_p_dout0;
            tmp_28_reg_1089 <= grp_fu_430_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state74)) begin
            pf_load_reg_1057 <= pf_q0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state69)) begin
            result_4_reg_1013 <= result_4_fu_529_p2;
            val_reg_1007 <= val_fu_522_p3;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state67)) begin
            select_ln18_2_reg_976 <= select_ln18_2_fu_341_p3;
            tmp_24_reg_971 <= add_ln486_1_fu_317_p2[32'd11];
            trunc_ln505_1_reg_966 <= trunc_ln505_1_fu_309_p1;
            xs_sign_1_reg_961 <= data_4_fu_287_p1[32'd63];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state68)) begin
            select_ln18_reg_996 <= select_ln18_fu_403_p3;
            tmp_22_reg_991 <= add_ln486_fu_379_p2[32'd11];
            trunc_ln505_reg_986 <= trunc_ln505_fu_371_p1;
            val_1_reg_1001 <= val_1_fu_463_p3;
            xs_sign_reg_981 <= data_fu_349_p1[32'd63];
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            tmp_25_reg_956 <= grp_fu_438_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            trunc_ln234_2_reg_1052 <= trunc_ln234_2_fu_705_p1;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state9)) begin
            xRay_2_reg_942 <= grp_fu_179_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state8)) begin
            yRay_2_reg_936 <= grp_fu_179_p_dout0;
        end
    end

    assign ap_ST_fsm_state10_blk = 1'b0;

    assign ap_ST_fsm_state11_blk = 1'b0;

    assign ap_ST_fsm_state12_blk = 1'b0;

    assign ap_ST_fsm_state13_blk = 1'b0;

    assign ap_ST_fsm_state14_blk = 1'b0;

    assign ap_ST_fsm_state15_blk = 1'b0;

    assign ap_ST_fsm_state16_blk = 1'b0;

    assign ap_ST_fsm_state17_blk = 1'b0;

    assign ap_ST_fsm_state18_blk = 1'b0;

    assign ap_ST_fsm_state19_blk = 1'b0;

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state20_blk = 1'b0;

    assign ap_ST_fsm_state21_blk = 1'b0;

    assign ap_ST_fsm_state22_blk = 1'b0;

    assign ap_ST_fsm_state23_blk = 1'b0;

    assign ap_ST_fsm_state24_blk = 1'b0;

    assign ap_ST_fsm_state25_blk = 1'b0;

    assign ap_ST_fsm_state26_blk = 1'b0;

    assign ap_ST_fsm_state27_blk = 1'b0;

    assign ap_ST_fsm_state28_blk = 1'b0;

    assign ap_ST_fsm_state29_blk = 1'b0;

    assign ap_ST_fsm_state2_blk  = 1'b0;

    assign ap_ST_fsm_state30_blk = 1'b0;

    assign ap_ST_fsm_state31_blk = 1'b0;

    assign ap_ST_fsm_state32_blk = 1'b0;

    assign ap_ST_fsm_state33_blk = 1'b0;

    assign ap_ST_fsm_state34_blk = 1'b0;

    assign ap_ST_fsm_state35_blk = 1'b0;

    assign ap_ST_fsm_state36_blk = 1'b0;

    assign ap_ST_fsm_state37_blk = 1'b0;

    assign ap_ST_fsm_state38_blk = 1'b0;

    assign ap_ST_fsm_state39_blk = 1'b0;

    assign ap_ST_fsm_state3_blk  = 1'b0;

    assign ap_ST_fsm_state40_blk = 1'b0;

    assign ap_ST_fsm_state41_blk = 1'b0;

    assign ap_ST_fsm_state42_blk = 1'b0;

    assign ap_ST_fsm_state43_blk = 1'b0;

    assign ap_ST_fsm_state44_blk = 1'b0;

    assign ap_ST_fsm_state45_blk = 1'b0;

    assign ap_ST_fsm_state46_blk = 1'b0;

    assign ap_ST_fsm_state47_blk = 1'b0;

    assign ap_ST_fsm_state48_blk = 1'b0;

    assign ap_ST_fsm_state49_blk = 1'b0;

    assign ap_ST_fsm_state4_blk  = 1'b0;

    assign ap_ST_fsm_state50_blk = 1'b0;

    assign ap_ST_fsm_state51_blk = 1'b0;

    assign ap_ST_fsm_state52_blk = 1'b0;

    assign ap_ST_fsm_state53_blk = 1'b0;

    assign ap_ST_fsm_state54_blk = 1'b0;

    assign ap_ST_fsm_state55_blk = 1'b0;

    assign ap_ST_fsm_state56_blk = 1'b0;

    assign ap_ST_fsm_state57_blk = 1'b0;

    assign ap_ST_fsm_state58_blk = 1'b0;

    assign ap_ST_fsm_state59_blk = 1'b0;

    assign ap_ST_fsm_state5_blk  = 1'b0;

    assign ap_ST_fsm_state60_blk = 1'b0;

    assign ap_ST_fsm_state61_blk = 1'b0;

    assign ap_ST_fsm_state62_blk = 1'b0;

    assign ap_ST_fsm_state63_blk = 1'b0;

    assign ap_ST_fsm_state64_blk = 1'b0;

    assign ap_ST_fsm_state65_blk = 1'b0;

    assign ap_ST_fsm_state66_blk = 1'b0;

    assign ap_ST_fsm_state67_blk = 1'b0;

    assign ap_ST_fsm_state68_blk = 1'b0;

    assign ap_ST_fsm_state69_blk = 1'b0;

    assign ap_ST_fsm_state6_blk  = 1'b0;

    assign ap_ST_fsm_state70_blk = 1'b0;

    assign ap_ST_fsm_state71_blk = 1'b0;

    assign ap_ST_fsm_state72_blk = 1'b0;

    assign ap_ST_fsm_state73_blk = 1'b0;

    assign ap_ST_fsm_state74_blk = 1'b0;

    assign ap_ST_fsm_state75_blk = 1'b0;

    assign ap_ST_fsm_state76_blk = 1'b0;

    assign ap_ST_fsm_state77_blk = 1'b0;

    assign ap_ST_fsm_state78_blk = 1'b0;

    assign ap_ST_fsm_state79_blk = 1'b0;

    assign ap_ST_fsm_state7_blk  = 1'b0;

    assign ap_ST_fsm_state80_blk = 1'b0;

    assign ap_ST_fsm_state81_blk = 1'b0;

    assign ap_ST_fsm_state82_blk = 1'b0;

    assign ap_ST_fsm_state8_blk  = 1'b0;

    assign ap_ST_fsm_state9_blk  = 1'b0;

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state81) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state81)) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_state82) | ((or_ln230_2_reg_1018 == 1'd0) & (1'b1 == ap_CS_fsm_state81)))) begin
            dist_1_out_ap_vld = 1'b1;
        end else begin
            dist_1_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_238_p0 = dist_fu_132;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_fu_238_p0 = xRay_1_fu_140;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_fu_238_p0 = yRay_1_fu_136;
        end else begin
            grp_fu_238_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            grp_fu_238_p1 = step;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_fu_238_p1 = xStep;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            grp_fu_238_p1 = yStep;
        end else begin
            grp_fu_238_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_fu_242_p0 = xRay_2_reg_942;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            grp_fu_242_p0 = yRay_2_reg_936;
        end else begin
            grp_fu_242_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state78)) begin
            grp_fu_246_p0 = occ_reg_1083;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_246_p0 = dist_1_reg_948;
        end else begin
            grp_fu_246_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state78)) begin
            grp_fu_246_p1 = bitcast_ln235;
        end else if ((1'b1 == ap_CS_fsm_state11)) begin
            grp_fu_246_p1 = empty;
        end else begin
            grp_fu_246_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state73)) begin
            pf_ce0 = 1'b1;
        end else begin
            pf_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
            ap_ST_fsm_state5: begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end
            ap_ST_fsm_state6: begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end
            ap_ST_fsm_state7: begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
            ap_ST_fsm_state8: begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
            ap_ST_fsm_state9: begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
            ap_ST_fsm_state10: begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
            ap_ST_fsm_state11: begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end
            ap_ST_fsm_state12: begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
            ap_ST_fsm_state13: begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
            ap_ST_fsm_state14: begin
                ap_NS_fsm = ap_ST_fsm_state15;
            end
            ap_ST_fsm_state15: begin
                ap_NS_fsm = ap_ST_fsm_state16;
            end
            ap_ST_fsm_state16: begin
                ap_NS_fsm = ap_ST_fsm_state17;
            end
            ap_ST_fsm_state17: begin
                ap_NS_fsm = ap_ST_fsm_state18;
            end
            ap_ST_fsm_state18: begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
            ap_ST_fsm_state19: begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
            ap_ST_fsm_state20: begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end
            ap_ST_fsm_state21: begin
                ap_NS_fsm = ap_ST_fsm_state22;
            end
            ap_ST_fsm_state22: begin
                ap_NS_fsm = ap_ST_fsm_state23;
            end
            ap_ST_fsm_state23: begin
                ap_NS_fsm = ap_ST_fsm_state24;
            end
            ap_ST_fsm_state24: begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end
            ap_ST_fsm_state25: begin
                ap_NS_fsm = ap_ST_fsm_state26;
            end
            ap_ST_fsm_state26: begin
                ap_NS_fsm = ap_ST_fsm_state27;
            end
            ap_ST_fsm_state27: begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
            ap_ST_fsm_state28: begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
            ap_ST_fsm_state29: begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end
            ap_ST_fsm_state30: begin
                ap_NS_fsm = ap_ST_fsm_state31;
            end
            ap_ST_fsm_state31: begin
                ap_NS_fsm = ap_ST_fsm_state32;
            end
            ap_ST_fsm_state32: begin
                ap_NS_fsm = ap_ST_fsm_state33;
            end
            ap_ST_fsm_state33: begin
                ap_NS_fsm = ap_ST_fsm_state34;
            end
            ap_ST_fsm_state34: begin
                ap_NS_fsm = ap_ST_fsm_state35;
            end
            ap_ST_fsm_state35: begin
                ap_NS_fsm = ap_ST_fsm_state36;
            end
            ap_ST_fsm_state36: begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
            ap_ST_fsm_state37: begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
            ap_ST_fsm_state38: begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end
            ap_ST_fsm_state39: begin
                ap_NS_fsm = ap_ST_fsm_state40;
            end
            ap_ST_fsm_state40: begin
                ap_NS_fsm = ap_ST_fsm_state41;
            end
            ap_ST_fsm_state41: begin
                ap_NS_fsm = ap_ST_fsm_state42;
            end
            ap_ST_fsm_state42: begin
                ap_NS_fsm = ap_ST_fsm_state43;
            end
            ap_ST_fsm_state43: begin
                ap_NS_fsm = ap_ST_fsm_state44;
            end
            ap_ST_fsm_state44: begin
                ap_NS_fsm = ap_ST_fsm_state45;
            end
            ap_ST_fsm_state45: begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
            ap_ST_fsm_state46: begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end
            ap_ST_fsm_state47: begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
            ap_ST_fsm_state48: begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
            ap_ST_fsm_state49: begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end
            ap_ST_fsm_state50: begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
            ap_ST_fsm_state51: begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end
            ap_ST_fsm_state52: begin
                ap_NS_fsm = ap_ST_fsm_state53;
            end
            ap_ST_fsm_state53: begin
                ap_NS_fsm = ap_ST_fsm_state54;
            end
            ap_ST_fsm_state54: begin
                ap_NS_fsm = ap_ST_fsm_state55;
            end
            ap_ST_fsm_state55: begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
            ap_ST_fsm_state56: begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
            ap_ST_fsm_state57: begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end
            ap_ST_fsm_state58: begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
            ap_ST_fsm_state59: begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end
            ap_ST_fsm_state60: begin
                ap_NS_fsm = ap_ST_fsm_state61;
            end
            ap_ST_fsm_state61: begin
                ap_NS_fsm = ap_ST_fsm_state62;
            end
            ap_ST_fsm_state62: begin
                ap_NS_fsm = ap_ST_fsm_state63;
            end
            ap_ST_fsm_state63: begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
            ap_ST_fsm_state64: begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end
            ap_ST_fsm_state65: begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
            ap_ST_fsm_state66: begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end
            ap_ST_fsm_state67: begin
                ap_NS_fsm = ap_ST_fsm_state68;
            end
            ap_ST_fsm_state68: begin
                ap_NS_fsm = ap_ST_fsm_state69;
            end
            ap_ST_fsm_state69: begin
                ap_NS_fsm = ap_ST_fsm_state70;
            end
            ap_ST_fsm_state70: begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
            ap_ST_fsm_state71: begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
            ap_ST_fsm_state72: begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end
            ap_ST_fsm_state73: begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
            ap_ST_fsm_state74: begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end
            ap_ST_fsm_state75: begin
                ap_NS_fsm = ap_ST_fsm_state76;
            end
            ap_ST_fsm_state76: begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end
            ap_ST_fsm_state77: begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end
            ap_ST_fsm_state78: begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
            ap_ST_fsm_state79: begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end
            ap_ST_fsm_state80: begin
                if (((or_ln235_3_fu_817_p2 == 1'd0) & (or_ln230_2_reg_1018 == 1'd0) & (1'b1 == ap_CS_fsm_state80))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else if (((or_ln230_2_reg_1018 == 1'd1) & (1'b1 == ap_CS_fsm_state80))) begin
                    ap_NS_fsm = ap_ST_fsm_state82;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state81;
                end
            end
            ap_ST_fsm_state81: begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
            ap_ST_fsm_state82: begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln234_fu_681_p2 = (zext_ln234_1_fu_677_p1 + 15'd16000);

    assign add_ln486_1_fu_317_p2 = ($signed(zext_ln486_1_fu_313_p1) + $signed(12'd3073));

    assign add_ln486_fu_379_p2 = ($signed(zext_ln486_fu_375_p1) + $signed(12'd3073));

    assign and_ln230_1_fu_595_p2 = (tmp_25_reg_956 & and_ln230_fu_589_p2);

    assign and_ln230_fu_589_p2 = (or_ln230_fu_579_p2 & or_ln230_1_fu_585_p2);

    assign and_ln235_1_fu_796_p2 = (or_ln235_2_fu_792_p2 & or_ln235_1_fu_788_p2);

    assign and_ln235_2_fu_802_p2 = (grp_fu_438_p_dout0 & and_ln235_1_fu_796_p2);

    assign and_ln235_fu_812_p2 = (tmp_28_reg_1089 & or_ln235_fu_808_p2);

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

    assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];

    assign ap_CS_fsm_state68 = ap_CS_fsm[32'd67];

    assign ap_CS_fsm_state69 = ap_CS_fsm[32'd68];

    assign ap_CS_fsm_state70 = ap_CS_fsm[32'd69];

    assign ap_CS_fsm_state72 = ap_CS_fsm[32'd71];

    assign ap_CS_fsm_state73 = ap_CS_fsm[32'd72];

    assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];

    assign ap_CS_fsm_state75 = ap_CS_fsm[32'd74];

    assign ap_CS_fsm_state77 = ap_CS_fsm[32'd76];

    assign ap_CS_fsm_state78 = ap_CS_fsm[32'd77];

    assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

    assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

    assign ap_CS_fsm_state81 = ap_CS_fsm[32'd80];

    assign ap_CS_fsm_state82 = ap_CS_fsm[32'd81];

    assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

    assign bitcast_ln230_fu_550_p1 = dist_1_reg_948;

    assign bitcast_ln234_fu_754_p1 = trunc_ln234_3_reg_1062;

    assign bitcast_ln235_1_fu_759_p1 = occ_reg_1083;

    assign data_4_fu_287_p1 = grp_fu_434_p_dout0;

    assign data_fu_349_p1 = grp_fu_434_p_dout0;

    assign dist_1_out = dist_1_reg_948;

    assign grp_fu_179_p_ce = 1'b1;

    assign grp_fu_179_p_din0 = grp_fu_238_p0;

    assign grp_fu_179_p_din1 = grp_fu_238_p1;

    assign grp_fu_179_p_opcode = 2'd0;

    assign grp_fu_427_p_ce = 1'b1;

    assign grp_fu_427_p_din0 = bitcast_ln234_fu_754_p1;

    assign grp_fu_430_p_ce = 1'b1;

    assign grp_fu_430_p_din0 = bitcast_ln234_fu_754_p1;

    assign grp_fu_430_p_din1 = 32'd3212836864;

    assign grp_fu_430_p_opcode = 5'd1;

    assign grp_fu_434_p_ce = 1'b1;

    assign grp_fu_434_p_din0 = grp_fu_242_p0;

    assign grp_fu_434_p_din1 = step;

    assign grp_fu_438_p_ce = 1'b1;

    assign grp_fu_438_p_din0 = grp_fu_246_p0;

    assign grp_fu_438_p_din1 = grp_fu_246_p1;

    assign grp_fu_438_p_opcode = 5'd3;

    assign grp_fu_834_p0 = grp_fu_834_p00;

    assign grp_fu_834_p00 = trunc_ln234_fu_638_p1;

    assign grp_fu_834_p1 = 22'd3200;

    assign grp_fu_834_p2 = grp_fu_834_p20;

    assign grp_fu_834_p20 = add_ln234_fu_681_p2;

    assign icmp_ln230_1_fu_567_p2 = ((tmp_s_fu_553_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln230_2_fu_614_p2 = ((result_fu_539_p3 > 32'd799) ? 1'b1 : 1'b0);

    assign icmp_ln230_3_fu_573_p2 = ((trunc_ln230_fu_563_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln230_4_fu_269_p2 = ((tmp_30 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln230_5_fu_274_p2 = ((trunc_ln230_1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln230_fu_600_p2 = (($signed(result_6_fu_545_p3) > $signed(32'd799)) ? 1'b1 : 1'b0);

    assign icmp_ln235_1_fu_748_p2 = ((trunc_ln235_fu_738_p1 == 23'd0) ? 1'b1 : 1'b0);

    assign icmp_ln235_2_fu_776_p2 = ((tmp_29_fu_762_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln235_3_fu_782_p2 = ((trunc_ln235_1_fu_772_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln235_4_fu_659_p2 = ((tmp_31_fu_650_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln235_5_fu_665_p2 = ((trunc_ln235_3 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln235_fu_742_p2 = ((tmp_27_fu_728_p4 != 8'd255) ? 1'b1 : 1'b0);

    assign lshr_ln18_1_fu_431_p2 = zext_ln15_1_fu_420_p1 >> zext_ln18_1_fu_427_p1;

    assign lshr_ln18_fu_490_p2 = zext_ln15_fu_479_p1 >> zext_ln18_fu_486_p1;

    assign lshr_ln234_1_fu_691_p4 = {{grp_fu_834_p3[21:5]}};

    assign lshr_ln234_fu_719_p2 = pf_load_reg_1057 >> zext_ln234_4_fu_715_p1;

    assign mantissa_1_fu_411_p4 = {{{{1'd1}, {trunc_ln505_1_reg_966}}}, {1'd0}};

    assign mantissa_fu_470_p4 = {{{{1'd1}, {trunc_ln505_reg_986}}}, {1'd0}};

    assign or_ln230_1_fu_585_p2 = (icmp_ln230_5_reg_921 | icmp_ln230_4_reg_916);

    assign or_ln230_2_fu_632_p2 = (or_ln230_4_fu_620_p2 | or_ln230_3_fu_626_p2);

    assign or_ln230_3_fu_626_p2 = (tmp_26_fu_606_p3 | icmp_ln230_2_fu_614_p2);

    assign or_ln230_4_fu_620_p2 = (icmp_ln230_fu_600_p2 | and_ln230_1_fu_595_p2);

    assign or_ln230_fu_579_p2 = (icmp_ln230_3_fu_573_p2 | icmp_ln230_1_fu_567_p2);

    assign or_ln235_1_fu_788_p2 = (icmp_ln235_3_reg_1099 | icmp_ln235_2_reg_1094);

    assign or_ln235_2_fu_792_p2 = (icmp_ln235_5_reg_1037 | icmp_ln235_4_reg_1032);

    assign or_ln235_3_fu_817_p2 = (and_ln235_fu_812_p2 | and_ln235_2_reg_1104);

    assign or_ln235_fu_808_p2 = (icmp_ln235_reg_1067 | icmp_ln235_1_reg_1072);

    assign pf_address0 = zext_ln234_3_fu_700_p1;

    assign result_1_fu_534_p2 = (32'd0 - val_reg_1007);

    assign result_4_fu_529_p2 = (32'd0 - val_1_reg_1001);

    assign result_6_fu_545_p3 = ((xs_sign_1_reg_961[0:0] == 1'b1) ? result_4_reg_1013 : val_1_reg_1001);

    assign result_fu_539_p3 = ((xs_sign_reg_981[0:0] == 1'b1) ? result_1_fu_534_p2 : val_reg_1007);

    assign select_ln18_2_fu_341_p3 = ((tmp_24_fu_323_p3[0:0] == 1'b1) ? sext_ln18_2_fu_337_p1 : add_ln486_1_fu_317_p2);

    assign select_ln18_fu_403_p3 = ((tmp_22_fu_385_p3[0:0] == 1'b1) ? sext_ln18_fu_399_p1 : add_ln486_fu_379_p2);

    assign sext_ln18_1_fu_483_p1 = $signed(select_ln18_reg_996);

    assign sext_ln18_2_fu_337_p1 = $signed(sub_ln18_1_fu_331_p2);

    assign sext_ln18_3_fu_424_p1 = $signed(select_ln18_2_reg_976);

    assign sext_ln18_fu_399_p1 = $signed(sub_ln18_fu_393_p2);

    assign shl_ln18_1_fu_437_p2 = zext_ln15_1_fu_420_p1 << zext_ln18_1_fu_427_p1;

    assign shl_ln18_fu_496_p2 = zext_ln15_fu_479_p1 << zext_ln18_fu_486_p1;

    assign shl_ln234_1_fu_708_p3 = {{trunc_ln234_2_reg_1052}, {3'd0}};

    assign shl_ln_fu_670_p3 = {{trunc_ln234_1_reg_1027}, {2'd0}};

    assign sub_ln18_1_fu_331_p2 = (11'd1023 - xs_exp_1_fu_299_p4);

    assign sub_ln18_fu_393_p2 = (11'd1023 - xs_exp_fu_361_p4);

    assign tmp_14_fu_502_p4 = {{lshr_ln18_fu_490_p2[84:53]}};

    assign tmp_15_fu_512_p4 = {{shl_ln18_fu_496_p2[84:53]}};

    assign tmp_16_fu_443_p4 = {{lshr_ln18_1_fu_431_p2[84:53]}};

    assign tmp_17_fu_453_p4 = {{shl_ln18_1_fu_437_p2[84:53]}};

    assign tmp_22_fu_385_p3 = add_ln486_fu_379_p2[32'd11];

    assign tmp_24_fu_323_p3 = add_ln486_1_fu_317_p2[32'd11];

    assign tmp_26_fu_606_p3 = result_6_fu_545_p3[32'd31];

    assign tmp_27_fu_728_p4 = {{lshr_ln234_fu_719_p2[30:23]}};

    assign tmp_29_fu_762_p4 = {{bitcast_ln235_1_fu_759_p1[62:52]}};

    assign tmp_31_fu_650_p4 = {{pf_load_6[190:180]}};

    assign tmp_s_fu_553_p4 = {{bitcast_ln230_fu_550_p1[62:52]}};

    assign trunc_ln230_fu_563_p1 = bitcast_ln230_fu_550_p1[51:0];

    assign trunc_ln234_1_fu_646_p1 = result_6_fu_545_p3[9:0];

    assign trunc_ln234_2_fu_705_p1 = grp_fu_834_p3[4:0];

    assign trunc_ln234_3_fu_724_p1 = lshr_ln234_fu_719_p2[31:0];

    assign trunc_ln234_fu_638_p1 = result_fu_539_p3[9:0];

    assign trunc_ln235_1_fu_772_p1 = bitcast_ln235_1_fu_759_p1[51:0];

    assign trunc_ln235_fu_738_p1 = lshr_ln234_fu_719_p2[22:0];

    assign trunc_ln505_1_fu_309_p1 = data_4_fu_287_p1[51:0];

    assign trunc_ln505_fu_371_p1 = data_fu_349_p1[51:0];

    assign val_1_fu_463_p3 = ((tmp_24_reg_971[0:0] == 1'b1) ? tmp_16_fu_443_p4 : tmp_17_fu_453_p4);

    assign val_fu_522_p3 = ((tmp_22_reg_991[0:0] == 1'b1) ? tmp_14_fu_502_p4 : tmp_15_fu_512_p4);

    assign xs_exp_1_fu_299_p4 = {{data_4_fu_287_p1[62:52]}};

    assign xs_exp_fu_361_p4 = {{data_fu_349_p1[62:52]}};

    assign zext_ln15_1_fu_420_p1 = mantissa_1_fu_411_p4;

    assign zext_ln15_fu_479_p1 = mantissa_fu_470_p4;

    assign zext_ln18_1_fu_427_p1 = $unsigned(sext_ln18_3_fu_424_p1);

    assign zext_ln18_fu_486_p1 = $unsigned(sext_ln18_1_fu_483_p1);

    assign zext_ln234_1_fu_677_p1 = shl_ln_fu_670_p3;

    assign zext_ln234_3_fu_700_p1 = lshr_ln234_1_fu_691_p4;

    assign zext_ln234_4_fu_715_p1 = shl_ln234_1_fu_708_p3;

    assign zext_ln486_1_fu_313_p1 = xs_exp_1_fu_299_p4;

    assign zext_ln486_fu_375_p1 = xs_exp_fu_361_p4;

endmodule  //main_rayCast_Pipeline_VITIS_LOOP_222_1
