/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_rpyxyzToH_double_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    x,
    y,
    z,
    H_0_0_address0,
    H_0_0_ce0,
    H_0_0_we0,
    H_0_0_d0,
    H_0_1_address0,
    H_0_1_ce0,
    H_0_1_we0,
    H_0_1_d0,
    H_0_2_address0,
    H_0_2_ce0,
    H_0_2_we0,
    H_0_2_d0,
    H_0_3_address0,
    H_0_3_ce0,
    H_0_3_we0,
    H_0_3_d0,
    H_1_0_address0,
    H_1_0_ce0,
    H_1_0_we0,
    H_1_0_d0,
    H_1_1_address0,
    H_1_1_ce0,
    H_1_1_we0,
    H_1_1_d0,
    H_1_2_address0,
    H_1_2_ce0,
    H_1_2_we0,
    H_1_2_d0,
    H_1_3_address0,
    H_1_3_ce0,
    H_1_3_we0,
    H_1_3_d0,
    H_2_0_address0,
    H_2_0_ce0,
    H_2_0_we0,
    H_2_0_d0,
    H_2_1_address0,
    H_2_1_ce0,
    H_2_1_we0,
    H_2_1_d0,
    H_2_2_address0,
    H_2_2_ce0,
    H_2_2_we0,
    H_2_2_d0,
    H_2_3_address0,
    H_2_3_ce0,
    H_2_3_we0,
    H_2_3_d0,
    H_3_0_address0,
    H_3_0_ce0,
    H_3_0_we0,
    H_3_0_d0,
    H_3_1_address0,
    H_3_1_ce0,
    H_3_1_we0,
    H_3_1_d0,
    H_3_2_address0,
    H_3_2_ce0,
    H_3_2_we0,
    H_3_2_d0,
    H_3_3_address0,
    H_3_3_ce0,
    H_3_3_we0,
    H_3_3_d0,
    H_offset
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] x;
    input [63:0] y;
    input [63:0] z;
    output [2:0] H_0_0_address0;
    output H_0_0_ce0;
    output H_0_0_we0;
    output [63:0] H_0_0_d0;
    output [2:0] H_0_1_address0;
    output H_0_1_ce0;
    output H_0_1_we0;
    output [63:0] H_0_1_d0;
    output [2:0] H_0_2_address0;
    output H_0_2_ce0;
    output H_0_2_we0;
    output [63:0] H_0_2_d0;
    output [2:0] H_0_3_address0;
    output H_0_3_ce0;
    output H_0_3_we0;
    output [63:0] H_0_3_d0;
    output [2:0] H_1_0_address0;
    output H_1_0_ce0;
    output H_1_0_we0;
    output [63:0] H_1_0_d0;
    output [2:0] H_1_1_address0;
    output H_1_1_ce0;
    output H_1_1_we0;
    output [63:0] H_1_1_d0;
    output [2:0] H_1_2_address0;
    output H_1_2_ce0;
    output H_1_2_we0;
    output [63:0] H_1_2_d0;
    output [2:0] H_1_3_address0;
    output H_1_3_ce0;
    output H_1_3_we0;
    output [63:0] H_1_3_d0;
    output [2:0] H_2_0_address0;
    output H_2_0_ce0;
    output H_2_0_we0;
    output [63:0] H_2_0_d0;
    output [2:0] H_2_1_address0;
    output H_2_1_ce0;
    output H_2_1_we0;
    output [63:0] H_2_1_d0;
    output [2:0] H_2_2_address0;
    output H_2_2_ce0;
    output H_2_2_we0;
    output [63:0] H_2_2_d0;
    output [2:0] H_2_3_address0;
    output H_2_3_ce0;
    output H_2_3_we0;
    output [63:0] H_2_3_d0;
    output [2:0] H_3_0_address0;
    output H_3_0_ce0;
    output H_3_0_we0;
    output [63:0] H_3_0_d0;
    output [2:0] H_3_1_address0;
    output H_3_1_ce0;
    output H_3_1_we0;
    output [63:0] H_3_1_d0;
    output [2:0] H_3_2_address0;
    output H_3_2_ce0;
    output H_3_2_we0;
    output [63:0] H_3_2_d0;
    output [2:0] H_3_3_address0;
    output H_3_3_ce0;
    output H_3_3_we0;
    output [63:0] H_3_3_d0;
    input [2:0] H_offset;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg H_0_0_ce0;
    reg H_0_0_we0;
    reg H_0_1_ce0;
    reg H_0_1_we0;
    reg H_0_2_ce0;
    reg H_0_2_we0;
    reg H_0_3_ce0;
    reg H_0_3_we0;
    reg H_1_0_ce0;
    reg H_1_0_we0;
    reg H_1_1_ce0;
    reg H_1_1_we0;
    reg H_1_2_ce0;
    reg H_1_2_we0;
    reg H_1_3_ce0;
    reg H_1_3_we0;
    reg H_2_0_ce0;
    reg H_2_0_we0;
    reg H_2_1_ce0;
    reg H_2_1_we0;
    reg H_2_2_ce0;
    reg H_2_2_we0;
    reg H_2_3_ce0;
    reg H_2_3_we0;
    reg H_3_0_ce0;
    reg H_3_0_we0;
    reg H_3_1_ce0;
    reg H_3_1_we0;
    reg H_3_2_ce0;
    reg H_3_2_we0;
    reg H_3_3_ce0;
    reg H_3_3_we0;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_enable_reg_pp0_iter27;
    reg    ap_enable_reg_pp0_iter28;
    reg    ap_enable_reg_pp0_iter29;
    reg    ap_enable_reg_pp0_iter30;
    reg    ap_enable_reg_pp0_iter31;
    reg    ap_enable_reg_pp0_iter32;
    reg    ap_enable_reg_pp0_iter33;
    reg    ap_enable_reg_pp0_iter34;
    reg    ap_enable_reg_pp0_iter35;
    reg    ap_enable_reg_pp0_iter36;
    reg    ap_enable_reg_pp0_iter37;
    reg    ap_enable_reg_pp0_iter38;
    reg    ap_enable_reg_pp0_iter39;
    reg    ap_enable_reg_pp0_iter40;
    reg    ap_enable_reg_pp0_iter41;
    reg    ap_enable_reg_pp0_iter42;
    reg    ap_enable_reg_pp0_iter43;
    reg    ap_enable_reg_pp0_iter44;
    reg    ap_enable_reg_pp0_iter45;
    reg    ap_enable_reg_pp0_iter46;
    reg    ap_enable_reg_pp0_iter47;
    reg    ap_enable_reg_pp0_iter48;
    reg    ap_enable_reg_pp0_iter49;
    reg    ap_enable_reg_pp0_iter50;
    reg    ap_enable_reg_pp0_iter51;
    reg    ap_enable_reg_pp0_iter52;
    reg    ap_enable_reg_pp0_iter53;
    reg    ap_enable_reg_pp0_iter54;
    reg    ap_enable_reg_pp0_iter55;
    reg    ap_enable_reg_pp0_iter56;
    reg    ap_enable_reg_pp0_iter57;
    reg    ap_enable_reg_pp0_iter58;
    reg    ap_enable_reg_pp0_iter59;
    reg    ap_enable_reg_pp0_iter60;
    reg    ap_enable_reg_pp0_iter61;
    reg    ap_enable_reg_pp0_iter62;
    reg    ap_enable_reg_pp0_iter63;
    reg    ap_enable_reg_pp0_iter64;
    reg    ap_enable_reg_pp0_iter65;
    reg    ap_enable_reg_pp0_iter66;
    reg    ap_enable_reg_pp0_iter67;
    reg    ap_enable_reg_pp0_iter68;
    reg    ap_enable_reg_pp0_iter69;
    reg    ap_enable_reg_pp0_iter70;
    reg    ap_enable_reg_pp0_iter71;
    reg    ap_enable_reg_pp0_iter72;
    reg    ap_enable_reg_pp0_iter73;
    reg    ap_enable_reg_pp0_iter74;
    reg    ap_enable_reg_pp0_iter75;
    reg    ap_enable_reg_pp0_iter76;
    reg    ap_enable_reg_pp0_iter77;
    reg    ap_idle_pp0;
    wire    ap_block_pp0_stage0_subdone;
    reg   [63:0] z_read_reg_820;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] z_read_reg_820_pp0_iter1_reg;
    reg   [63:0] z_read_reg_820_pp0_iter2_reg;
    reg   [63:0] z_read_reg_820_pp0_iter3_reg;
    reg   [63:0] z_read_reg_820_pp0_iter4_reg;
    reg   [63:0] z_read_reg_820_pp0_iter5_reg;
    reg   [63:0] z_read_reg_820_pp0_iter6_reg;
    reg   [63:0] z_read_reg_820_pp0_iter7_reg;
    reg   [63:0] z_read_reg_820_pp0_iter8_reg;
    reg   [63:0] z_read_reg_820_pp0_iter9_reg;
    reg   [63:0] z_read_reg_820_pp0_iter10_reg;
    reg   [63:0] z_read_reg_820_pp0_iter11_reg;
    reg   [63:0] z_read_reg_820_pp0_iter12_reg;
    reg   [63:0] z_read_reg_820_pp0_iter13_reg;
    reg   [63:0] z_read_reg_820_pp0_iter14_reg;
    reg   [63:0] z_read_reg_820_pp0_iter15_reg;
    reg   [63:0] z_read_reg_820_pp0_iter16_reg;
    reg   [63:0] z_read_reg_820_pp0_iter17_reg;
    reg   [63:0] z_read_reg_820_pp0_iter18_reg;
    reg   [63:0] z_read_reg_820_pp0_iter19_reg;
    reg   [63:0] z_read_reg_820_pp0_iter20_reg;
    reg   [63:0] y_read_reg_826;
    reg   [63:0] y_read_reg_826_pp0_iter1_reg;
    reg   [63:0] y_read_reg_826_pp0_iter2_reg;
    reg   [63:0] y_read_reg_826_pp0_iter3_reg;
    reg   [63:0] y_read_reg_826_pp0_iter4_reg;
    reg   [63:0] y_read_reg_826_pp0_iter5_reg;
    reg   [63:0] y_read_reg_826_pp0_iter6_reg;
    reg   [63:0] y_read_reg_826_pp0_iter7_reg;
    reg   [63:0] y_read_reg_826_pp0_iter8_reg;
    reg   [63:0] y_read_reg_826_pp0_iter9_reg;
    reg   [63:0] y_read_reg_826_pp0_iter10_reg;
    reg   [63:0] y_read_reg_826_pp0_iter11_reg;
    reg   [63:0] y_read_reg_826_pp0_iter12_reg;
    reg   [63:0] y_read_reg_826_pp0_iter13_reg;
    reg   [63:0] y_read_reg_826_pp0_iter14_reg;
    reg   [63:0] y_read_reg_826_pp0_iter15_reg;
    reg   [63:0] y_read_reg_826_pp0_iter16_reg;
    reg   [63:0] y_read_reg_826_pp0_iter17_reg;
    reg   [63:0] y_read_reg_826_pp0_iter18_reg;
    reg   [63:0] y_read_reg_826_pp0_iter19_reg;
    reg   [63:0] y_read_reg_826_pp0_iter20_reg;
    reg   [63:0] x_read_reg_832;
    reg   [63:0] x_read_reg_832_pp0_iter1_reg;
    reg   [63:0] x_read_reg_832_pp0_iter2_reg;
    reg   [63:0] x_read_reg_832_pp0_iter3_reg;
    reg   [63:0] x_read_reg_832_pp0_iter4_reg;
    reg   [63:0] x_read_reg_832_pp0_iter5_reg;
    reg   [63:0] x_read_reg_832_pp0_iter6_reg;
    reg   [63:0] x_read_reg_832_pp0_iter7_reg;
    reg   [63:0] x_read_reg_832_pp0_iter8_reg;
    reg   [63:0] x_read_reg_832_pp0_iter9_reg;
    reg   [63:0] x_read_reg_832_pp0_iter10_reg;
    reg   [63:0] x_read_reg_832_pp0_iter11_reg;
    reg   [63:0] x_read_reg_832_pp0_iter12_reg;
    reg   [63:0] x_read_reg_832_pp0_iter13_reg;
    reg   [63:0] x_read_reg_832_pp0_iter14_reg;
    reg   [63:0] x_read_reg_832_pp0_iter15_reg;
    reg   [63:0] x_read_reg_832_pp0_iter16_reg;
    reg   [63:0] x_read_reg_832_pp0_iter17_reg;
    reg   [63:0] x_read_reg_832_pp0_iter18_reg;
    reg   [63:0] x_read_reg_832_pp0_iter19_reg;
    reg   [63:0] x_read_reg_832_pp0_iter20_reg;
    wire   [63:0] H_offset_cast_fu_812_p1;
    reg   [63:0] H_offset_cast_reg_838;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter1_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter2_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter3_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter4_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter5_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter6_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter7_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter8_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter9_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter10_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter11_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter12_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter13_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter14_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter15_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter16_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter17_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter18_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter19_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter20_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter21_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter22_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter23_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter24_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter25_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter26_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter27_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter28_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter29_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter30_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter31_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter32_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter33_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter34_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter35_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter36_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter37_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter38_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter39_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter40_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter41_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter42_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter43_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter44_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter45_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter46_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter47_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter48_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter49_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter50_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter51_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter52_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter53_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter54_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter55_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter56_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter57_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter58_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter59_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter60_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter61_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter62_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter63_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter64_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter65_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter66_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter67_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter68_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter69_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter70_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter71_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter72_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter73_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter74_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter75_reg;
    reg   [63:0] H_offset_cast_reg_838_pp0_iter76_reg;
    wire   [63:0] grp_fu_659_p2;
    reg   [63:0] mul_i_0_0_3_reg_854;
    wire   [63:0] grp_fu_665_p2;
    reg   [63:0] mul_i_1_0_3_reg_860;
    wire   [63:0] grp_fu_671_p2;
    reg   [63:0] mul_i_2_0_3_reg_866;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter7_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter8_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter9_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter10_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter11_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter12_reg;
    reg   [63:0] mul_i_2_0_3_reg_866_pp0_iter13_reg;
    wire   [63:0] grp_fu_288_p2;
    reg   [63:0] add_i_0_0_3_reg_872;
    wire   [63:0] grp_fu_293_p2;
    reg   [63:0] add_i_0_1_3_reg_878;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter14_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter15_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter16_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter17_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter18_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter19_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter20_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter21_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter22_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter23_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter24_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter25_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter26_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter27_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter28_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter29_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter30_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter31_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter32_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter33_reg;
    reg   [63:0] add_i_0_1_3_reg_878_pp0_iter34_reg;
    wire   [63:0] grp_fu_298_p2;
    reg   [63:0] add_i_1_0_3_reg_886;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter14_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter15_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter16_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter17_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter18_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter19_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter20_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter21_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter22_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter23_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter24_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter25_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter26_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter27_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter28_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter29_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter30_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter31_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter32_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter33_reg;
    reg   [63:0] add_i_1_0_3_reg_886_pp0_iter34_reg;
    wire   [63:0] grp_fu_303_p2;
    reg   [63:0] add_i_1_1_3_reg_894;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter14_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter15_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter16_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter17_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter18_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter19_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter20_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter21_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter22_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter23_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter24_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter25_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter26_reg;
    reg   [63:0] add_i_1_1_3_reg_894_pp0_iter27_reg;
    wire   [63:0] grp_fu_308_p2;
    reg   [63:0] add_i_2_0_3_reg_900;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter14_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter15_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter16_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter17_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter18_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter19_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter20_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter21_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter22_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter23_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter24_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter25_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter26_reg;
    reg   [63:0] add_i_2_0_3_reg_900_pp0_iter27_reg;
    wire   [63:0] grp_fu_313_p2;
    reg   [63:0] add_i_2_2_3_reg_907;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter21_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter22_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter23_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter24_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter25_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter26_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter27_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter28_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter29_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter30_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter31_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter32_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter33_reg;
    reg   [63:0] add_i_2_2_3_reg_907_pp0_iter34_reg;
    wire   [63:0] grp_fu_318_p2;
    reg   [63:0] add_i1_reg_914;
    wire   [63:0] grp_fu_677_p2;
    reg   [63:0] mul_i1_0_0_1_reg_919;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter21_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter22_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter23_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter24_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter25_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter26_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter27_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter28_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter29_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter30_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter31_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter32_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter33_reg;
    reg   [63:0] mul_i1_0_0_1_reg_919_pp0_iter34_reg;
    wire   [63:0] grp_fu_682_p2;
    reg   [63:0] mul_i1_0_1_reg_927;
    wire   [63:0] grp_fu_687_p2;
    reg   [63:0] mul_i1_1_0_1_reg_932;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter21_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter22_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter23_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter24_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter25_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter26_reg;
    reg   [63:0] mul_i1_1_0_1_reg_932_pp0_iter27_reg;
    wire   [63:0] grp_fu_692_p2;
    reg   [63:0] mul_i1_1_1_reg_938;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter21_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter22_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter23_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter24_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter25_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter26_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter27_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter28_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter29_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter30_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter31_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter32_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter33_reg;
    reg   [63:0] mul_i1_1_1_reg_938_pp0_iter34_reg;
    wire   [63:0] grp_fu_697_p2;
    reg   [63:0] mul_i1_2_0_1_reg_945;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter21_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter22_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter23_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter24_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter25_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter26_reg;
    reg   [63:0] mul_i1_2_0_1_reg_945_pp0_iter27_reg;
    wire   [63:0] grp_fu_323_p2;
    reg   [63:0] add_i_0_3_3_reg_952;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter28_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter29_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter30_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter31_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter32_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter33_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter34_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter35_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter36_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter37_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter38_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter39_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter40_reg;
    reg   [63:0] add_i_0_3_3_reg_952_pp0_iter41_reg;
    wire   [63:0] grp_fu_328_p2;
    reg   [63:0] add_i_1_3_3_reg_958;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter28_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter29_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter30_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter31_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter32_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter33_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter34_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter35_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter36_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter37_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter38_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter39_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter40_reg;
    reg   [63:0] add_i_1_3_3_reg_958_pp0_iter41_reg;
    wire   [63:0] grp_fu_333_p2;
    reg   [63:0] add_i_2_3_3_reg_964;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter28_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter29_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter30_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter31_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter32_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter33_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter34_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter35_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter36_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter37_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter38_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter39_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter40_reg;
    reg   [63:0] add_i_2_3_3_reg_964_pp0_iter41_reg;
    wire   [63:0] grp_fu_338_p2;
    reg   [63:0] add_i1_0_0_1_reg_970;
    wire   [63:0] grp_fu_702_p2;
    reg   [63:0] mul_i1_0_0_2_reg_975;
    wire   [63:0] grp_fu_342_p2;
    reg   [63:0] add_i1_0_1_reg_980;
    wire   [63:0] grp_fu_347_p2;
    reg   [63:0] add_i1_1_0_1_reg_986;
    wire   [63:0] grp_fu_707_p2;
    reg   [63:0] mul_i1_1_0_2_reg_991;
    wire   [63:0] grp_fu_351_p2;
    reg   [63:0] add_i1_1_1_reg_996;
    wire   [63:0] grp_fu_356_p2;
    reg   [63:0] add_i1_2_0_1_reg_1002;
    wire   [63:0] grp_fu_712_p2;
    reg   [63:0] mul_i1_2_0_2_reg_1007;
    wire   [63:0] grp_fu_360_p2;
    reg   [63:0] add_i1_2_1_reg_1012;
    wire   [63:0] grp_fu_365_p2;
    reg   [63:0] add_i1_0_0_2_reg_1018;
    wire   [63:0] grp_fu_717_p2;
    reg   [63:0] mul_i1_0_0_3_reg_1023;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter35_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter36_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter37_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter38_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter39_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter40_reg;
    reg   [63:0] mul_i1_0_0_3_reg_1023_pp0_iter41_reg;
    wire   [63:0] grp_fu_369_p2;
    reg   [63:0] add_i1_0_1_1_reg_1030;
    wire   [63:0] grp_fu_373_p2;
    reg   [63:0] add_i1_0_2_1_reg_1035;
    wire   [63:0] grp_fu_377_p2;
    reg   [63:0] add_i1_1_0_2_reg_1041;
    wire   [63:0] grp_fu_722_p2;
    reg   [63:0] mul_i1_1_0_3_reg_1046;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter35_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter36_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter37_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter38_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter39_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter40_reg;
    reg   [63:0] mul_i1_1_0_3_reg_1046_pp0_iter41_reg;
    wire   [63:0] grp_fu_381_p2;
    reg   [63:0] add_i1_1_1_1_reg_1053;
    wire   [63:0] grp_fu_385_p2;
    reg   [63:0] add_i1_1_2_1_reg_1058;
    wire   [63:0] grp_fu_389_p2;
    reg   [63:0] add_i1_2_0_2_reg_1064;
    wire   [63:0] grp_fu_727_p2;
    reg   [63:0] mul_i1_2_0_3_reg_1069;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter35_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter36_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter37_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter38_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter39_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter40_reg;
    reg   [63:0] mul_i1_2_0_3_reg_1069_pp0_iter41_reg;
    wire   [63:0] grp_fu_393_p2;
    reg   [63:0] add_i1_2_1_1_reg_1076;
    wire   [63:0] grp_fu_732_p2;
    reg   [63:0] mul_i1_2_1_2_reg_1081;
    wire   [63:0] grp_fu_397_p2;
    reg   [63:0] add_i1_2_2_1_reg_1087;
    wire   [63:0] grp_fu_401_p2;
    reg   [63:0] add_i1_0_0_3_reg_1093;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter42_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter43_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter44_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter45_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter46_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter47_reg;
    reg   [63:0] add_i1_0_0_3_reg_1093_pp0_iter48_reg;
    wire   [63:0] grp_fu_405_p2;
    reg   [63:0] add_i1_0_1_2_reg_1099;
    wire   [63:0] grp_fu_409_p2;
    reg   [63:0] add_i1_0_2_2_reg_1104;
    wire   [63:0] grp_fu_413_p2;
    reg   [63:0] add_i1_0_3_2_reg_1109;
    wire   [63:0] grp_fu_417_p2;
    reg   [63:0] add_i1_1_0_3_reg_1114;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter42_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter43_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter44_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter45_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter46_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter47_reg;
    reg   [63:0] add_i1_1_0_3_reg_1114_pp0_iter48_reg;
    wire   [63:0] grp_fu_421_p2;
    reg   [63:0] add_i1_1_1_2_reg_1120;
    wire   [63:0] grp_fu_425_p2;
    reg   [63:0] add_i1_1_2_2_reg_1125;
    wire   [63:0] grp_fu_429_p2;
    reg   [63:0] add_i1_1_3_2_reg_1130;
    wire   [63:0] grp_fu_433_p2;
    reg   [63:0] add_i1_2_0_3_reg_1135;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter42_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter43_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter44_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter45_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter46_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter47_reg;
    reg   [63:0] add_i1_2_0_3_reg_1135_pp0_iter48_reg;
    wire   [63:0] grp_fu_437_p2;
    reg   [63:0] add_i1_2_1_2_reg_1141;
    wire   [63:0] grp_fu_441_p2;
    reg   [63:0] add_i1_2_2_2_reg_1146;
    wire   [63:0] grp_fu_445_p2;
    reg   [63:0] add_i1_2_3_2_reg_1151;
    wire   [63:0] grp_fu_449_p2;
    reg   [63:0] add_i1_0_1_3_reg_1156;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter49_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter50_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter51_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter52_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter53_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter54_reg;
    reg   [63:0] add_i1_0_1_3_reg_1156_pp0_iter55_reg;
    wire   [63:0] grp_fu_453_p2;
    reg   [63:0] add_i1_0_2_3_reg_1163;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter49_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter50_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter51_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter52_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter53_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter54_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter55_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter56_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter57_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter58_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter59_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter60_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter61_reg;
    reg   [63:0] add_i1_0_2_3_reg_1163_pp0_iter62_reg;
    wire   [63:0] grp_fu_457_p2;
    reg   [63:0] add_i1_0_3_3_reg_1169;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter49_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter50_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter51_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter52_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter53_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter54_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter55_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter56_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter57_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter58_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter59_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter60_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter61_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter62_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter63_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter64_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter65_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter66_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter67_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter68_reg;
    reg   [63:0] add_i1_0_3_3_reg_1169_pp0_iter69_reg;
    wire   [63:0] grp_fu_461_p2;
    reg   [63:0] add_i1_1_1_3_reg_1175;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter49_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter50_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter51_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter52_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter53_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter54_reg;
    reg   [63:0] add_i1_1_1_3_reg_1175_pp0_iter55_reg;
    wire   [63:0] grp_fu_465_p2;
    reg   [63:0] add_i1_1_2_3_reg_1182;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter49_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter50_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter51_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter52_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter53_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter54_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter55_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter56_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter57_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter58_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter59_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter60_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter61_reg;
    reg   [63:0] add_i1_1_2_3_reg_1182_pp0_iter62_reg;
    wire   [63:0] grp_fu_469_p2;
    reg   [63:0] add_i1_1_3_3_reg_1188;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter49_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter50_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter51_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter52_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter53_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter54_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter55_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter56_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter57_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter58_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter59_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter60_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter61_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter62_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter63_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter64_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter65_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter66_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter67_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter68_reg;
    reg   [63:0] add_i1_1_3_3_reg_1188_pp0_iter69_reg;
    wire   [63:0] grp_fu_473_p2;
    reg   [63:0] add_i1_2_1_3_reg_1194;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter49_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter50_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter51_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter52_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter53_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter54_reg;
    reg   [63:0] add_i1_2_1_3_reg_1194_pp0_iter55_reg;
    wire   [63:0] grp_fu_477_p2;
    reg   [63:0] add_i1_2_2_3_reg_1201;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter49_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter50_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter51_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter52_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter53_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter54_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter55_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter56_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter57_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter58_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter59_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter60_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter61_reg;
    reg   [63:0] add_i1_2_2_3_reg_1201_pp0_iter62_reg;
    wire   [63:0] grp_fu_481_p2;
    reg   [63:0] add_i1_2_3_3_reg_1207;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter49_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter50_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter51_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter52_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter53_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter54_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter55_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter56_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter57_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter58_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter59_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter60_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter61_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter62_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter63_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter64_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter65_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter66_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter67_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter68_reg;
    reg   [63:0] add_i1_2_3_3_reg_1207_pp0_iter69_reg;
    wire   [63:0] grp_fu_737_p2;
    reg   [63:0] mul_i2_0_1_reg_1213;
    wire   [63:0] grp_fu_742_p2;
    reg   [63:0] mul_i2_1_1_reg_1218;
    wire   [63:0] grp_fu_747_p2;
    reg   [63:0] mul_i2_2_1_reg_1223;
    wire   [63:0] grp_fu_485_p2;
    reg   [63:0] add_i2_reg_1228;
    wire   [63:0] grp_fu_752_p2;
    reg   [63:0] mul_i2_0_0_1_reg_1233;
    wire   [63:0] grp_fu_490_p2;
    reg   [63:0] add_i2_0_1_reg_1239;
    wire   [63:0] grp_fu_757_p2;
    reg   [63:0] mul_i2_0_2_1_reg_1246;
    wire   [63:0] grp_fu_495_p2;
    reg   [63:0] add_i2_1_reg_1251;
    wire   [63:0] grp_fu_762_p2;
    reg   [63:0] mul_i2_1_0_1_reg_1256;
    wire   [63:0] grp_fu_500_p2;
    reg   [63:0] add_i2_1_1_reg_1262;
    wire   [63:0] grp_fu_767_p2;
    reg   [63:0] mul_i2_1_2_1_reg_1269;
    wire   [63:0] grp_fu_505_p2;
    reg   [63:0] add_i2_2_reg_1274;
    wire   [63:0] grp_fu_772_p2;
    reg   [63:0] mul_i2_2_0_1_reg_1279;
    wire   [63:0] grp_fu_510_p2;
    reg   [63:0] add_i2_2_1_reg_1285;
    wire   [63:0] grp_fu_777_p2;
    reg   [63:0] mul_i2_2_2_1_reg_1292;
    wire   [63:0] grp_fu_515_p2;
    reg   [63:0] add_i2_0_0_1_reg_1297;
    wire   [63:0] grp_fu_782_p2;
    reg   [63:0] mul_i2_0_0_2_reg_1302;
    wire   [63:0] grp_fu_519_p2;
    reg   [63:0] add_i2_0_1_1_reg_1309;
    wire   [63:0] grp_fu_523_p2;
    reg   [63:0] add_i2_0_2_1_reg_1314;
    wire   [63:0] grp_fu_527_p2;
    reg   [63:0] add_i2_0_3_1_reg_1319;
    wire   [63:0] grp_fu_531_p2;
    reg   [63:0] add_i2_1_0_1_reg_1324;
    wire   [63:0] grp_fu_787_p2;
    reg   [63:0] mul_i2_1_0_2_reg_1329;
    wire   [63:0] grp_fu_535_p2;
    reg   [63:0] add_i2_1_1_1_reg_1336;
    wire   [63:0] grp_fu_539_p2;
    reg   [63:0] add_i2_1_2_1_reg_1341;
    wire   [63:0] grp_fu_543_p2;
    reg   [63:0] add_i2_1_3_1_reg_1346;
    wire   [63:0] grp_fu_547_p2;
    reg   [63:0] add_i2_2_0_1_reg_1351;
    wire   [63:0] grp_fu_792_p2;
    reg   [63:0] mul_i2_2_0_2_reg_1356;
    wire   [63:0] grp_fu_551_p2;
    reg   [63:0] add_i2_2_1_1_reg_1363;
    wire   [63:0] grp_fu_555_p2;
    reg   [63:0] add_i2_2_2_1_reg_1368;
    wire   [63:0] grp_fu_559_p2;
    reg   [63:0] add_i2_2_3_1_reg_1373;
    wire   [63:0] grp_fu_563_p2;
    reg   [63:0] add_i2_0_0_2_reg_1378;
    wire   [63:0] grp_fu_797_p2;
    reg   [63:0] mul_i2_0_0_3_reg_1383;
    wire   [63:0] grp_fu_567_p2;
    reg   [63:0] add_i2_0_1_2_reg_1390;
    wire   [63:0] grp_fu_571_p2;
    reg   [63:0] add_i2_0_2_2_reg_1395;
    wire   [63:0] grp_fu_575_p2;
    reg   [63:0] add_i2_0_3_2_reg_1400;
    wire   [63:0] grp_fu_579_p2;
    reg   [63:0] add_i2_1_0_2_reg_1405;
    wire   [63:0] grp_fu_802_p2;
    reg   [63:0] mul_i2_1_0_3_reg_1410;
    wire   [63:0] grp_fu_583_p2;
    reg   [63:0] add_i2_1_1_2_reg_1417;
    wire   [63:0] grp_fu_587_p2;
    reg   [63:0] add_i2_1_2_2_reg_1422;
    wire   [63:0] grp_fu_591_p2;
    reg   [63:0] add_i2_1_3_2_reg_1427;
    wire   [63:0] grp_fu_595_p2;
    reg   [63:0] add_i2_2_0_2_reg_1432;
    wire   [63:0] grp_fu_807_p2;
    reg   [63:0] mul_i2_2_0_3_reg_1437;
    wire   [63:0] grp_fu_599_p2;
    reg   [63:0] add_i2_2_1_2_reg_1444;
    wire   [63:0] grp_fu_603_p2;
    reg   [63:0] add_i2_2_2_2_reg_1449;
    wire   [63:0] grp_fu_607_p2;
    reg   [63:0] add_i2_2_3_2_reg_1454;
    wire   [63:0] grp_fu_611_p2;
    reg   [63:0] add_i2_0_0_3_reg_1459;
    wire   [63:0] grp_fu_615_p2;
    reg   [63:0] add_i2_0_1_3_reg_1464;
    wire   [63:0] grp_fu_619_p2;
    reg   [63:0] add_i2_0_2_3_reg_1469;
    wire   [63:0] grp_fu_623_p2;
    reg   [63:0] add_i2_0_3_3_reg_1474;
    wire   [63:0] grp_fu_627_p2;
    reg   [63:0] add_i2_1_0_3_reg_1479;
    wire   [63:0] grp_fu_631_p2;
    reg   [63:0] add_i2_1_1_3_reg_1484;
    wire   [63:0] grp_fu_635_p2;
    reg   [63:0] add_i2_1_2_3_reg_1489;
    wire   [63:0] grp_fu_639_p2;
    reg   [63:0] add_i2_1_3_3_reg_1494;
    wire   [63:0] grp_fu_643_p2;
    reg   [63:0] add_i2_2_0_3_reg_1499;
    wire   [63:0] grp_fu_647_p2;
    reg   [63:0] add_i2_2_1_3_reg_1504;
    wire   [63:0] grp_fu_651_p2;
    reg   [63:0] add_i2_2_2_3_reg_1509;
    wire   [63:0] grp_fu_655_p2;
    reg   [63:0] add_i2_2_3_3_reg_1514;
    wire    ap_block_pp0_stage0;
    reg   [0:0] ap_NS_fsm;
    reg    ap_idle_pp0_0to76;
    reg    ap_reset_idle_pp0;
    wire    ap_enable_pp0;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter27 = 1'b0;
        #0 ap_enable_reg_pp0_iter28 = 1'b0;
        #0 ap_enable_reg_pp0_iter29 = 1'b0;
        #0 ap_enable_reg_pp0_iter30 = 1'b0;
        #0 ap_enable_reg_pp0_iter31 = 1'b0;
        #0 ap_enable_reg_pp0_iter32 = 1'b0;
        #0 ap_enable_reg_pp0_iter33 = 1'b0;
        #0 ap_enable_reg_pp0_iter34 = 1'b0;
        #0 ap_enable_reg_pp0_iter35 = 1'b0;
        #0 ap_enable_reg_pp0_iter36 = 1'b0;
        #0 ap_enable_reg_pp0_iter37 = 1'b0;
        #0 ap_enable_reg_pp0_iter38 = 1'b0;
        #0 ap_enable_reg_pp0_iter39 = 1'b0;
        #0 ap_enable_reg_pp0_iter40 = 1'b0;
        #0 ap_enable_reg_pp0_iter41 = 1'b0;
        #0 ap_enable_reg_pp0_iter42 = 1'b0;
        #0 ap_enable_reg_pp0_iter43 = 1'b0;
        #0 ap_enable_reg_pp0_iter44 = 1'b0;
        #0 ap_enable_reg_pp0_iter45 = 1'b0;
        #0 ap_enable_reg_pp0_iter46 = 1'b0;
        #0 ap_enable_reg_pp0_iter47 = 1'b0;
        #0 ap_enable_reg_pp0_iter48 = 1'b0;
        #0 ap_enable_reg_pp0_iter49 = 1'b0;
        #0 ap_enable_reg_pp0_iter50 = 1'b0;
        #0 ap_enable_reg_pp0_iter51 = 1'b0;
        #0 ap_enable_reg_pp0_iter52 = 1'b0;
        #0 ap_enable_reg_pp0_iter53 = 1'b0;
        #0 ap_enable_reg_pp0_iter54 = 1'b0;
        #0 ap_enable_reg_pp0_iter55 = 1'b0;
        #0 ap_enable_reg_pp0_iter56 = 1'b0;
        #0 ap_enable_reg_pp0_iter57 = 1'b0;
        #0 ap_enable_reg_pp0_iter58 = 1'b0;
        #0 ap_enable_reg_pp0_iter59 = 1'b0;
        #0 ap_enable_reg_pp0_iter60 = 1'b0;
        #0 ap_enable_reg_pp0_iter61 = 1'b0;
        #0 ap_enable_reg_pp0_iter62 = 1'b0;
        #0 ap_enable_reg_pp0_iter63 = 1'b0;
        #0 ap_enable_reg_pp0_iter64 = 1'b0;
        #0 ap_enable_reg_pp0_iter65 = 1'b0;
        #0 ap_enable_reg_pp0_iter66 = 1'b0;
        #0 ap_enable_reg_pp0_iter67 = 1'b0;
        #0 ap_enable_reg_pp0_iter68 = 1'b0;
        #0 ap_enable_reg_pp0_iter69 = 1'b0;
        #0 ap_enable_reg_pp0_iter70 = 1'b0;
        #0 ap_enable_reg_pp0_iter71 = 1'b0;
        #0 ap_enable_reg_pp0_iter72 = 1'b0;
        #0 ap_enable_reg_pp0_iter73 = 1'b0;
        #0 ap_enable_reg_pp0_iter74 = 1'b0;
        #0 ap_enable_reg_pp0_iter75 = 1'b0;
        #0 ap_enable_reg_pp0_iter76 = 1'b0;
        #0 ap_enable_reg_pp0_iter77 = 1'b0;
    end

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U154 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_854),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_288_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U155 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_0_0_3_reg_854),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_293_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U156 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_1_0_3_reg_860),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_298_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U157 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_1_0_3_reg_860),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_303_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U158 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_2_0_3_reg_866),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_308_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U159 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i_2_0_3_reg_866_pp0_iter13_reg),
        .din1(64'd4607182418800017408),
        .ce(1'b1),
        .dout(grp_fu_313_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U160 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_872),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_318_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U161 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x_read_reg_832_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_323_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U162 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(y_read_reg_826_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_328_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U163 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(z_read_reg_820_pp0_iter20_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_333_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U164 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_reg_914),
        .din1(mul_i1_0_0_1_reg_919),
        .ce(1'b1),
        .dout(grp_fu_338_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U165 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_0_1_reg_927),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_342_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U166 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_886_pp0_iter20_reg),
        .din1(mul_i1_1_0_1_reg_932),
        .ce(1'b1),
        .dout(grp_fu_347_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U167 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_1_1_reg_938),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_351_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U168 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_0_3_reg_900_pp0_iter20_reg),
        .din1(mul_i1_2_0_1_reg_945),
        .ce(1'b1),
        .dout(grp_fu_356_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U169 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i1_2_0_1_reg_945),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_360_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U170 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_1_reg_970),
        .din1(mul_i1_0_0_2_reg_975),
        .ce(1'b1),
        .dout(grp_fu_365_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U171 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_980),
        .din1(add_i_0_1_3_reg_878_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_369_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U172 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_reg_980),
        .din1(mul_i1_0_0_1_reg_919_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_373_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U173 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_1_reg_986),
        .din1(mul_i1_1_0_2_reg_991),
        .ce(1'b1),
        .dout(grp_fu_377_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U174 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_996),
        .din1(add_i_1_1_3_reg_894_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_381_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U175 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_reg_996),
        .din1(mul_i1_1_0_1_reg_932_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_385_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U176 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_1_reg_1002),
        .din1(mul_i1_2_0_2_reg_1007),
        .ce(1'b1),
        .dout(grp_fu_389_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U177 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_reg_1012),
        .din1(add_i_2_0_3_reg_900_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_393_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U178 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_reg_1012),
        .din1(mul_i1_2_0_1_reg_945_pp0_iter27_reg),
        .ce(1'b1),
        .dout(grp_fu_397_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U179 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_2_reg_1018),
        .din1(mul_i1_0_0_3_reg_1023),
        .ce(1'b1),
        .dout(grp_fu_401_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U180 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_1_reg_1030),
        .din1(mul_i1_0_0_1_reg_919_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_405_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U181 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_1035),
        .din1(add_i_0_1_3_reg_878_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_409_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U182 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_1_reg_1035),
        .din1(mul_i1_0_0_1_reg_919_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_413_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U183 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_2_reg_1041),
        .din1(mul_i1_1_0_3_reg_1046),
        .ce(1'b1),
        .dout(grp_fu_417_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U184 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_1_reg_1053),
        .din1(mul_i1_1_1_reg_938_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_421_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U185 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_1058),
        .din1(add_i_1_0_3_reg_886_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_425_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U186 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_1_reg_1058),
        .din1(mul_i1_1_1_reg_938_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_429_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U187 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_2_reg_1064),
        .din1(mul_i1_2_0_3_reg_1069),
        .ce(1'b1),
        .dout(grp_fu_433_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U188 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_1_reg_1076),
        .din1(mul_i1_2_1_2_reg_1081),
        .ce(1'b1),
        .dout(grp_fu_437_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U189 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_1087),
        .din1(add_i_2_2_3_reg_907_pp0_iter34_reg),
        .ce(1'b1),
        .dout(grp_fu_441_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U190 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_1_reg_1087),
        .din1(mul_i1_2_1_2_reg_1081),
        .ce(1'b1),
        .dout(grp_fu_445_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U191 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_2_reg_1099),
        .din1(mul_i1_0_0_3_reg_1023_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_449_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U192 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_2_reg_1104),
        .din1(mul_i1_0_0_3_reg_1023_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_453_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U193 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_2_reg_1109),
        .din1(add_i_0_3_3_reg_952_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_457_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U194 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_2_reg_1120),
        .din1(mul_i1_1_0_3_reg_1046_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_461_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U195 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_2_reg_1125),
        .din1(mul_i1_1_0_3_reg_1046_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_465_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U196 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_2_reg_1130),
        .din1(add_i_1_3_3_reg_958_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_469_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U197 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_2_reg_1141),
        .din1(mul_i1_2_0_3_reg_1069_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_473_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U198 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_2_reg_1146),
        .din1(mul_i1_2_0_3_reg_1069_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_477_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U199 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_2_reg_1151),
        .din1(add_i_2_3_3_reg_964_pp0_iter41_reg),
        .ce(1'b1),
        .dout(grp_fu_481_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U200 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_1093_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_485_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U201 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_0_1_reg_1213),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_490_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U202 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_1114_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_495_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U203 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_1_1_reg_1218),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_500_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U204 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_1135_pp0_iter48_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_505_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U205 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(mul_i2_2_1_reg_1223),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_510_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U206 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_reg_1228),
        .din1(mul_i2_0_0_1_reg_1233),
        .ce(1'b1),
        .dout(grp_fu_515_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U207 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_1239),
        .din1(add_i1_0_1_3_reg_1156_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_519_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U208 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_1239),
        .din1(mul_i2_0_2_1_reg_1246),
        .ce(1'b1),
        .dout(grp_fu_523_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U209 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_reg_1239),
        .din1(mul_i2_0_0_1_reg_1233),
        .ce(1'b1),
        .dout(grp_fu_527_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U210 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_reg_1251),
        .din1(mul_i2_1_0_1_reg_1256),
        .ce(1'b1),
        .dout(grp_fu_531_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U211 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_1262),
        .din1(add_i1_1_1_3_reg_1175_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_535_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U212 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_1262),
        .din1(mul_i2_1_2_1_reg_1269),
        .ce(1'b1),
        .dout(grp_fu_539_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U213 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_reg_1262),
        .din1(mul_i2_1_0_1_reg_1256),
        .ce(1'b1),
        .dout(grp_fu_543_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U214 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_reg_1274),
        .din1(mul_i2_2_0_1_reg_1279),
        .ce(1'b1),
        .dout(grp_fu_547_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U215 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_1285),
        .din1(add_i1_2_1_3_reg_1194_pp0_iter55_reg),
        .ce(1'b1),
        .dout(grp_fu_551_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U216 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_1285),
        .din1(mul_i2_2_2_1_reg_1292),
        .ce(1'b1),
        .dout(grp_fu_555_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U217 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_reg_1285),
        .din1(mul_i2_2_0_1_reg_1279),
        .ce(1'b1),
        .dout(grp_fu_559_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U218 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_1_reg_1297),
        .din1(mul_i2_0_0_2_reg_1302),
        .ce(1'b1),
        .dout(grp_fu_563_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U219 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_1_reg_1309),
        .din1(mul_i2_0_0_2_reg_1302),
        .ce(1'b1),
        .dout(grp_fu_567_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U220 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_1_reg_1314),
        .din1(add_i1_0_2_3_reg_1163_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_571_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U221 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_1_reg_1319),
        .din1(mul_i2_0_0_2_reg_1302),
        .ce(1'b1),
        .dout(grp_fu_575_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U222 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_1_reg_1324),
        .din1(mul_i2_1_0_2_reg_1329),
        .ce(1'b1),
        .dout(grp_fu_579_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U223 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_1_reg_1336),
        .din1(mul_i2_1_0_2_reg_1329),
        .ce(1'b1),
        .dout(grp_fu_583_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U224 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_1_reg_1341),
        .din1(add_i1_1_2_3_reg_1182_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_587_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U225 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_1_reg_1346),
        .din1(mul_i2_1_0_2_reg_1329),
        .ce(1'b1),
        .dout(grp_fu_591_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U226 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_1_reg_1351),
        .din1(mul_i2_2_0_2_reg_1356),
        .ce(1'b1),
        .dout(grp_fu_595_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U227 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_1_reg_1363),
        .din1(mul_i2_2_0_2_reg_1356),
        .ce(1'b1),
        .dout(grp_fu_599_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U228 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_1_reg_1368),
        .din1(add_i1_2_2_3_reg_1201_pp0_iter62_reg),
        .ce(1'b1),
        .dout(grp_fu_603_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U229 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_1_reg_1373),
        .din1(mul_i2_2_0_2_reg_1356),
        .ce(1'b1),
        .dout(grp_fu_607_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U230 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_0_2_reg_1378),
        .din1(mul_i2_0_0_3_reg_1383),
        .ce(1'b1),
        .dout(grp_fu_611_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U231 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_1_2_reg_1390),
        .din1(mul_i2_0_0_3_reg_1383),
        .ce(1'b1),
        .dout(grp_fu_615_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U232 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_2_2_reg_1395),
        .din1(mul_i2_0_0_3_reg_1383),
        .ce(1'b1),
        .dout(grp_fu_619_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U233 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_0_3_2_reg_1400),
        .din1(add_i1_0_3_3_reg_1169_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_623_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U234 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_0_2_reg_1405),
        .din1(mul_i2_1_0_3_reg_1410),
        .ce(1'b1),
        .dout(grp_fu_627_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U235 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_1_2_reg_1417),
        .din1(mul_i2_1_0_3_reg_1410),
        .ce(1'b1),
        .dout(grp_fu_631_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U236 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_2_2_reg_1422),
        .din1(mul_i2_1_0_3_reg_1410),
        .ce(1'b1),
        .dout(grp_fu_635_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U237 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_1_3_2_reg_1427),
        .din1(add_i1_1_3_3_reg_1188_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_639_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U238 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_0_2_reg_1432),
        .din1(mul_i2_2_0_3_reg_1437),
        .ce(1'b1),
        .dout(grp_fu_643_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U239 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_1_2_reg_1444),
        .din1(mul_i2_2_0_3_reg_1437),
        .ce(1'b1),
        .dout(grp_fu_647_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U240 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_2_2_reg_1449),
        .din1(mul_i2_2_0_3_reg_1437),
        .ce(1'b1),
        .dout(grp_fu_651_p2)
    );

    main_dadd_64ns_64ns_64_7_full_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadd_64ns_64ns_64_7_full_dsp_1_U241 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i2_2_3_2_reg_1454),
        .din1(add_i1_2_3_3_reg_1207_pp0_iter69_reg),
        .ce(1'b1),
        .dout(grp_fu_655_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U242 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(x),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_659_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U243 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(y),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_665_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U244 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(z),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_671_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U245 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_878),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_677_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U246 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_0_3_reg_872),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_682_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U247 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_1_3_reg_894),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_687_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U248 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_886),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_692_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U249 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_0_3_reg_900),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_697_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U250 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_1_3_reg_878_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_702_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U251 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_0_3_reg_886_pp0_iter20_reg),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_707_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U252 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_2_3_reg_907),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_712_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U253 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_0_3_3_reg_952),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_717_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U254 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_1_3_3_reg_958),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_722_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U255 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_3_3_reg_964),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_727_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U256 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i_2_2_3_reg_907_pp0_iter27_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_732_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U257 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_0_3_reg_1093),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_737_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U258 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_0_3_reg_1114),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_742_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U259 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_0_3_reg_1135),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_747_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U260 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_1156),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_752_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U261 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_1_3_reg_1156),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_757_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U262 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_1175),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_762_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U263 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_1_3_reg_1175),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_767_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U264 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_1194),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_772_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U265 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_1_3_reg_1194),
        .din1(64'd9223372036854775808),
        .ce(1'b1),
        .dout(grp_fu_777_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U266 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_2_3_reg_1163_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_782_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U267 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_2_3_reg_1182_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_787_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U268 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_2_3_reg_1201_pp0_iter55_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_792_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U269 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_0_3_3_reg_1169_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_797_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U270 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_1_3_3_reg_1188_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_802_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U271 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_i1_2_3_3_reg_1207_pp0_iter62_reg),
        .din1(64'd0),
        .ce(1'b1),
        .dout(grp_fu_807_p2)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
                ap_enable_reg_pp0_iter1 <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter27 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter28 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter29 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter30 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter31 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter32 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter33 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter33 <= ap_enable_reg_pp0_iter32;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter34 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter34 <= ap_enable_reg_pp0_iter33;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter35 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter35 <= ap_enable_reg_pp0_iter34;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter36 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter36 <= ap_enable_reg_pp0_iter35;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter37 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter37 <= ap_enable_reg_pp0_iter36;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter38 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter38 <= ap_enable_reg_pp0_iter37;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter39 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter39 <= ap_enable_reg_pp0_iter38;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter40 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter40 <= ap_enable_reg_pp0_iter39;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter41 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter41 <= ap_enable_reg_pp0_iter40;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter42 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter42 <= ap_enable_reg_pp0_iter41;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter43 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter43 <= ap_enable_reg_pp0_iter42;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter44 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter44 <= ap_enable_reg_pp0_iter43;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter45 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter45 <= ap_enable_reg_pp0_iter44;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter46 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter46 <= ap_enable_reg_pp0_iter45;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter47 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter47 <= ap_enable_reg_pp0_iter46;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter48 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter48 <= ap_enable_reg_pp0_iter47;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter49 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter49 <= ap_enable_reg_pp0_iter48;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter50 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter50 <= ap_enable_reg_pp0_iter49;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter51 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter51 <= ap_enable_reg_pp0_iter50;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter52 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter52 <= ap_enable_reg_pp0_iter51;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter53 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter53 <= ap_enable_reg_pp0_iter52;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter54 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter54 <= ap_enable_reg_pp0_iter53;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter55 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter55 <= ap_enable_reg_pp0_iter54;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter56 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter56 <= ap_enable_reg_pp0_iter55;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter57 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter57 <= ap_enable_reg_pp0_iter56;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter58 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter58 <= ap_enable_reg_pp0_iter57;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter59 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter59 <= ap_enable_reg_pp0_iter58;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter60 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter60 <= ap_enable_reg_pp0_iter59;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter61 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter61 <= ap_enable_reg_pp0_iter60;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter62 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter62 <= ap_enable_reg_pp0_iter61;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter63 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter63 <= ap_enable_reg_pp0_iter62;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter64 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter64 <= ap_enable_reg_pp0_iter63;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter65 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter65 <= ap_enable_reg_pp0_iter64;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter66 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter66 <= ap_enable_reg_pp0_iter65;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter67 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter67 <= ap_enable_reg_pp0_iter66;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter68 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter68 <= ap_enable_reg_pp0_iter67;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter69 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter69 <= ap_enable_reg_pp0_iter68;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter70 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter70 <= ap_enable_reg_pp0_iter69;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter71 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter71 <= ap_enable_reg_pp0_iter70;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter72 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter72 <= ap_enable_reg_pp0_iter71;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter73 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter73 <= ap_enable_reg_pp0_iter72;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter74 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter74 <= ap_enable_reg_pp0_iter73;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter75 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter75 <= ap_enable_reg_pp0_iter74;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter76 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter76 <= ap_enable_reg_pp0_iter75;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter77 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter77 <= ap_enable_reg_pp0_iter76;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_offset_cast_reg_838[2 : 0] <= H_offset_cast_fu_812_p1[2 : 0];
            H_offset_cast_reg_838_pp0_iter1_reg[2 : 0] <= H_offset_cast_reg_838[2 : 0];
            x_read_reg_832 <= x;
            x_read_reg_832_pp0_iter1_reg <= x_read_reg_832;
            y_read_reg_826 <= y;
            y_read_reg_826_pp0_iter1_reg <= y_read_reg_826;
            z_read_reg_820 <= z;
            z_read_reg_820_pp0_iter1_reg <= z_read_reg_820;
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b0 == ap_block_pp0_stage0_11001)) begin
            H_offset_cast_reg_838_pp0_iter10_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter9_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter11_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter10_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter12_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter11_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter13_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter12_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter14_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter13_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter15_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter14_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter16_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter15_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter17_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter16_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter18_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter17_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter19_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter18_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter20_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter19_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter21_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter20_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter22_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter21_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter23_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter22_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter24_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter23_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter25_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter24_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter26_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter25_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter27_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter26_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter28_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter27_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter29_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter28_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter2_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter1_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter30_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter29_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter31_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter30_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter32_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter31_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter33_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter32_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter34_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter33_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter35_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter34_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter36_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter35_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter37_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter36_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter38_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter37_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter39_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter38_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter3_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter2_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter40_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter39_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter41_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter40_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter42_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter41_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter43_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter42_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter44_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter43_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter45_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter44_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter46_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter45_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter47_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter46_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter48_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter47_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter49_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter48_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter4_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter3_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter50_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter49_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter51_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter50_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter52_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter51_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter53_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter52_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter54_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter53_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter55_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter54_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter56_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter55_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter57_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter56_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter58_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter57_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter59_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter58_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter5_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter4_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter60_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter59_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter61_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter60_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter62_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter61_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter63_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter62_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter64_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter63_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter65_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter64_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter66_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter65_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter67_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter66_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter68_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter67_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter69_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter68_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter6_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter5_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter70_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter69_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter71_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter70_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter72_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter71_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter73_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter72_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter74_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter73_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter75_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter74_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter76_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter75_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter7_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter6_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter8_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter7_reg[2 : 0];
            H_offset_cast_reg_838_pp0_iter9_reg[2 : 0] <= H_offset_cast_reg_838_pp0_iter8_reg[2 : 0];
            add_i1_0_0_1_reg_970 <= grp_fu_338_p2;
            add_i1_0_0_2_reg_1018 <= grp_fu_365_p2;
            add_i1_0_0_3_reg_1093 <= grp_fu_401_p2;
            add_i1_0_0_3_reg_1093_pp0_iter42_reg <= add_i1_0_0_3_reg_1093;
            add_i1_0_0_3_reg_1093_pp0_iter43_reg <= add_i1_0_0_3_reg_1093_pp0_iter42_reg;
            add_i1_0_0_3_reg_1093_pp0_iter44_reg <= add_i1_0_0_3_reg_1093_pp0_iter43_reg;
            add_i1_0_0_3_reg_1093_pp0_iter45_reg <= add_i1_0_0_3_reg_1093_pp0_iter44_reg;
            add_i1_0_0_3_reg_1093_pp0_iter46_reg <= add_i1_0_0_3_reg_1093_pp0_iter45_reg;
            add_i1_0_0_3_reg_1093_pp0_iter47_reg <= add_i1_0_0_3_reg_1093_pp0_iter46_reg;
            add_i1_0_0_3_reg_1093_pp0_iter48_reg <= add_i1_0_0_3_reg_1093_pp0_iter47_reg;
            add_i1_0_1_1_reg_1030 <= grp_fu_369_p2;
            add_i1_0_1_2_reg_1099 <= grp_fu_405_p2;
            add_i1_0_1_3_reg_1156 <= grp_fu_449_p2;
            add_i1_0_1_3_reg_1156_pp0_iter49_reg <= add_i1_0_1_3_reg_1156;
            add_i1_0_1_3_reg_1156_pp0_iter50_reg <= add_i1_0_1_3_reg_1156_pp0_iter49_reg;
            add_i1_0_1_3_reg_1156_pp0_iter51_reg <= add_i1_0_1_3_reg_1156_pp0_iter50_reg;
            add_i1_0_1_3_reg_1156_pp0_iter52_reg <= add_i1_0_1_3_reg_1156_pp0_iter51_reg;
            add_i1_0_1_3_reg_1156_pp0_iter53_reg <= add_i1_0_1_3_reg_1156_pp0_iter52_reg;
            add_i1_0_1_3_reg_1156_pp0_iter54_reg <= add_i1_0_1_3_reg_1156_pp0_iter53_reg;
            add_i1_0_1_3_reg_1156_pp0_iter55_reg <= add_i1_0_1_3_reg_1156_pp0_iter54_reg;
            add_i1_0_1_reg_980 <= grp_fu_342_p2;
            add_i1_0_2_1_reg_1035 <= grp_fu_373_p2;
            add_i1_0_2_2_reg_1104 <= grp_fu_409_p2;
            add_i1_0_2_3_reg_1163 <= grp_fu_453_p2;
            add_i1_0_2_3_reg_1163_pp0_iter49_reg <= add_i1_0_2_3_reg_1163;
            add_i1_0_2_3_reg_1163_pp0_iter50_reg <= add_i1_0_2_3_reg_1163_pp0_iter49_reg;
            add_i1_0_2_3_reg_1163_pp0_iter51_reg <= add_i1_0_2_3_reg_1163_pp0_iter50_reg;
            add_i1_0_2_3_reg_1163_pp0_iter52_reg <= add_i1_0_2_3_reg_1163_pp0_iter51_reg;
            add_i1_0_2_3_reg_1163_pp0_iter53_reg <= add_i1_0_2_3_reg_1163_pp0_iter52_reg;
            add_i1_0_2_3_reg_1163_pp0_iter54_reg <= add_i1_0_2_3_reg_1163_pp0_iter53_reg;
            add_i1_0_2_3_reg_1163_pp0_iter55_reg <= add_i1_0_2_3_reg_1163_pp0_iter54_reg;
            add_i1_0_2_3_reg_1163_pp0_iter56_reg <= add_i1_0_2_3_reg_1163_pp0_iter55_reg;
            add_i1_0_2_3_reg_1163_pp0_iter57_reg <= add_i1_0_2_3_reg_1163_pp0_iter56_reg;
            add_i1_0_2_3_reg_1163_pp0_iter58_reg <= add_i1_0_2_3_reg_1163_pp0_iter57_reg;
            add_i1_0_2_3_reg_1163_pp0_iter59_reg <= add_i1_0_2_3_reg_1163_pp0_iter58_reg;
            add_i1_0_2_3_reg_1163_pp0_iter60_reg <= add_i1_0_2_3_reg_1163_pp0_iter59_reg;
            add_i1_0_2_3_reg_1163_pp0_iter61_reg <= add_i1_0_2_3_reg_1163_pp0_iter60_reg;
            add_i1_0_2_3_reg_1163_pp0_iter62_reg <= add_i1_0_2_3_reg_1163_pp0_iter61_reg;
            add_i1_0_3_2_reg_1109 <= grp_fu_413_p2;
            add_i1_0_3_3_reg_1169 <= grp_fu_457_p2;
            add_i1_0_3_3_reg_1169_pp0_iter49_reg <= add_i1_0_3_3_reg_1169;
            add_i1_0_3_3_reg_1169_pp0_iter50_reg <= add_i1_0_3_3_reg_1169_pp0_iter49_reg;
            add_i1_0_3_3_reg_1169_pp0_iter51_reg <= add_i1_0_3_3_reg_1169_pp0_iter50_reg;
            add_i1_0_3_3_reg_1169_pp0_iter52_reg <= add_i1_0_3_3_reg_1169_pp0_iter51_reg;
            add_i1_0_3_3_reg_1169_pp0_iter53_reg <= add_i1_0_3_3_reg_1169_pp0_iter52_reg;
            add_i1_0_3_3_reg_1169_pp0_iter54_reg <= add_i1_0_3_3_reg_1169_pp0_iter53_reg;
            add_i1_0_3_3_reg_1169_pp0_iter55_reg <= add_i1_0_3_3_reg_1169_pp0_iter54_reg;
            add_i1_0_3_3_reg_1169_pp0_iter56_reg <= add_i1_0_3_3_reg_1169_pp0_iter55_reg;
            add_i1_0_3_3_reg_1169_pp0_iter57_reg <= add_i1_0_3_3_reg_1169_pp0_iter56_reg;
            add_i1_0_3_3_reg_1169_pp0_iter58_reg <= add_i1_0_3_3_reg_1169_pp0_iter57_reg;
            add_i1_0_3_3_reg_1169_pp0_iter59_reg <= add_i1_0_3_3_reg_1169_pp0_iter58_reg;
            add_i1_0_3_3_reg_1169_pp0_iter60_reg <= add_i1_0_3_3_reg_1169_pp0_iter59_reg;
            add_i1_0_3_3_reg_1169_pp0_iter61_reg <= add_i1_0_3_3_reg_1169_pp0_iter60_reg;
            add_i1_0_3_3_reg_1169_pp0_iter62_reg <= add_i1_0_3_3_reg_1169_pp0_iter61_reg;
            add_i1_0_3_3_reg_1169_pp0_iter63_reg <= add_i1_0_3_3_reg_1169_pp0_iter62_reg;
            add_i1_0_3_3_reg_1169_pp0_iter64_reg <= add_i1_0_3_3_reg_1169_pp0_iter63_reg;
            add_i1_0_3_3_reg_1169_pp0_iter65_reg <= add_i1_0_3_3_reg_1169_pp0_iter64_reg;
            add_i1_0_3_3_reg_1169_pp0_iter66_reg <= add_i1_0_3_3_reg_1169_pp0_iter65_reg;
            add_i1_0_3_3_reg_1169_pp0_iter67_reg <= add_i1_0_3_3_reg_1169_pp0_iter66_reg;
            add_i1_0_3_3_reg_1169_pp0_iter68_reg <= add_i1_0_3_3_reg_1169_pp0_iter67_reg;
            add_i1_0_3_3_reg_1169_pp0_iter69_reg <= add_i1_0_3_3_reg_1169_pp0_iter68_reg;
            add_i1_1_0_1_reg_986 <= grp_fu_347_p2;
            add_i1_1_0_2_reg_1041 <= grp_fu_377_p2;
            add_i1_1_0_3_reg_1114 <= grp_fu_417_p2;
            add_i1_1_0_3_reg_1114_pp0_iter42_reg <= add_i1_1_0_3_reg_1114;
            add_i1_1_0_3_reg_1114_pp0_iter43_reg <= add_i1_1_0_3_reg_1114_pp0_iter42_reg;
            add_i1_1_0_3_reg_1114_pp0_iter44_reg <= add_i1_1_0_3_reg_1114_pp0_iter43_reg;
            add_i1_1_0_3_reg_1114_pp0_iter45_reg <= add_i1_1_0_3_reg_1114_pp0_iter44_reg;
            add_i1_1_0_3_reg_1114_pp0_iter46_reg <= add_i1_1_0_3_reg_1114_pp0_iter45_reg;
            add_i1_1_0_3_reg_1114_pp0_iter47_reg <= add_i1_1_0_3_reg_1114_pp0_iter46_reg;
            add_i1_1_0_3_reg_1114_pp0_iter48_reg <= add_i1_1_0_3_reg_1114_pp0_iter47_reg;
            add_i1_1_1_1_reg_1053 <= grp_fu_381_p2;
            add_i1_1_1_2_reg_1120 <= grp_fu_421_p2;
            add_i1_1_1_3_reg_1175 <= grp_fu_461_p2;
            add_i1_1_1_3_reg_1175_pp0_iter49_reg <= add_i1_1_1_3_reg_1175;
            add_i1_1_1_3_reg_1175_pp0_iter50_reg <= add_i1_1_1_3_reg_1175_pp0_iter49_reg;
            add_i1_1_1_3_reg_1175_pp0_iter51_reg <= add_i1_1_1_3_reg_1175_pp0_iter50_reg;
            add_i1_1_1_3_reg_1175_pp0_iter52_reg <= add_i1_1_1_3_reg_1175_pp0_iter51_reg;
            add_i1_1_1_3_reg_1175_pp0_iter53_reg <= add_i1_1_1_3_reg_1175_pp0_iter52_reg;
            add_i1_1_1_3_reg_1175_pp0_iter54_reg <= add_i1_1_1_3_reg_1175_pp0_iter53_reg;
            add_i1_1_1_3_reg_1175_pp0_iter55_reg <= add_i1_1_1_3_reg_1175_pp0_iter54_reg;
            add_i1_1_1_reg_996 <= grp_fu_351_p2;
            add_i1_1_2_1_reg_1058 <= grp_fu_385_p2;
            add_i1_1_2_2_reg_1125 <= grp_fu_425_p2;
            add_i1_1_2_3_reg_1182 <= grp_fu_465_p2;
            add_i1_1_2_3_reg_1182_pp0_iter49_reg <= add_i1_1_2_3_reg_1182;
            add_i1_1_2_3_reg_1182_pp0_iter50_reg <= add_i1_1_2_3_reg_1182_pp0_iter49_reg;
            add_i1_1_2_3_reg_1182_pp0_iter51_reg <= add_i1_1_2_3_reg_1182_pp0_iter50_reg;
            add_i1_1_2_3_reg_1182_pp0_iter52_reg <= add_i1_1_2_3_reg_1182_pp0_iter51_reg;
            add_i1_1_2_3_reg_1182_pp0_iter53_reg <= add_i1_1_2_3_reg_1182_pp0_iter52_reg;
            add_i1_1_2_3_reg_1182_pp0_iter54_reg <= add_i1_1_2_3_reg_1182_pp0_iter53_reg;
            add_i1_1_2_3_reg_1182_pp0_iter55_reg <= add_i1_1_2_3_reg_1182_pp0_iter54_reg;
            add_i1_1_2_3_reg_1182_pp0_iter56_reg <= add_i1_1_2_3_reg_1182_pp0_iter55_reg;
            add_i1_1_2_3_reg_1182_pp0_iter57_reg <= add_i1_1_2_3_reg_1182_pp0_iter56_reg;
            add_i1_1_2_3_reg_1182_pp0_iter58_reg <= add_i1_1_2_3_reg_1182_pp0_iter57_reg;
            add_i1_1_2_3_reg_1182_pp0_iter59_reg <= add_i1_1_2_3_reg_1182_pp0_iter58_reg;
            add_i1_1_2_3_reg_1182_pp0_iter60_reg <= add_i1_1_2_3_reg_1182_pp0_iter59_reg;
            add_i1_1_2_3_reg_1182_pp0_iter61_reg <= add_i1_1_2_3_reg_1182_pp0_iter60_reg;
            add_i1_1_2_3_reg_1182_pp0_iter62_reg <= add_i1_1_2_3_reg_1182_pp0_iter61_reg;
            add_i1_1_3_2_reg_1130 <= grp_fu_429_p2;
            add_i1_1_3_3_reg_1188 <= grp_fu_469_p2;
            add_i1_1_3_3_reg_1188_pp0_iter49_reg <= add_i1_1_3_3_reg_1188;
            add_i1_1_3_3_reg_1188_pp0_iter50_reg <= add_i1_1_3_3_reg_1188_pp0_iter49_reg;
            add_i1_1_3_3_reg_1188_pp0_iter51_reg <= add_i1_1_3_3_reg_1188_pp0_iter50_reg;
            add_i1_1_3_3_reg_1188_pp0_iter52_reg <= add_i1_1_3_3_reg_1188_pp0_iter51_reg;
            add_i1_1_3_3_reg_1188_pp0_iter53_reg <= add_i1_1_3_3_reg_1188_pp0_iter52_reg;
            add_i1_1_3_3_reg_1188_pp0_iter54_reg <= add_i1_1_3_3_reg_1188_pp0_iter53_reg;
            add_i1_1_3_3_reg_1188_pp0_iter55_reg <= add_i1_1_3_3_reg_1188_pp0_iter54_reg;
            add_i1_1_3_3_reg_1188_pp0_iter56_reg <= add_i1_1_3_3_reg_1188_pp0_iter55_reg;
            add_i1_1_3_3_reg_1188_pp0_iter57_reg <= add_i1_1_3_3_reg_1188_pp0_iter56_reg;
            add_i1_1_3_3_reg_1188_pp0_iter58_reg <= add_i1_1_3_3_reg_1188_pp0_iter57_reg;
            add_i1_1_3_3_reg_1188_pp0_iter59_reg <= add_i1_1_3_3_reg_1188_pp0_iter58_reg;
            add_i1_1_3_3_reg_1188_pp0_iter60_reg <= add_i1_1_3_3_reg_1188_pp0_iter59_reg;
            add_i1_1_3_3_reg_1188_pp0_iter61_reg <= add_i1_1_3_3_reg_1188_pp0_iter60_reg;
            add_i1_1_3_3_reg_1188_pp0_iter62_reg <= add_i1_1_3_3_reg_1188_pp0_iter61_reg;
            add_i1_1_3_3_reg_1188_pp0_iter63_reg <= add_i1_1_3_3_reg_1188_pp0_iter62_reg;
            add_i1_1_3_3_reg_1188_pp0_iter64_reg <= add_i1_1_3_3_reg_1188_pp0_iter63_reg;
            add_i1_1_3_3_reg_1188_pp0_iter65_reg <= add_i1_1_3_3_reg_1188_pp0_iter64_reg;
            add_i1_1_3_3_reg_1188_pp0_iter66_reg <= add_i1_1_3_3_reg_1188_pp0_iter65_reg;
            add_i1_1_3_3_reg_1188_pp0_iter67_reg <= add_i1_1_3_3_reg_1188_pp0_iter66_reg;
            add_i1_1_3_3_reg_1188_pp0_iter68_reg <= add_i1_1_3_3_reg_1188_pp0_iter67_reg;
            add_i1_1_3_3_reg_1188_pp0_iter69_reg <= add_i1_1_3_3_reg_1188_pp0_iter68_reg;
            add_i1_2_0_1_reg_1002 <= grp_fu_356_p2;
            add_i1_2_0_2_reg_1064 <= grp_fu_389_p2;
            add_i1_2_0_3_reg_1135 <= grp_fu_433_p2;
            add_i1_2_0_3_reg_1135_pp0_iter42_reg <= add_i1_2_0_3_reg_1135;
            add_i1_2_0_3_reg_1135_pp0_iter43_reg <= add_i1_2_0_3_reg_1135_pp0_iter42_reg;
            add_i1_2_0_3_reg_1135_pp0_iter44_reg <= add_i1_2_0_3_reg_1135_pp0_iter43_reg;
            add_i1_2_0_3_reg_1135_pp0_iter45_reg <= add_i1_2_0_3_reg_1135_pp0_iter44_reg;
            add_i1_2_0_3_reg_1135_pp0_iter46_reg <= add_i1_2_0_3_reg_1135_pp0_iter45_reg;
            add_i1_2_0_3_reg_1135_pp0_iter47_reg <= add_i1_2_0_3_reg_1135_pp0_iter46_reg;
            add_i1_2_0_3_reg_1135_pp0_iter48_reg <= add_i1_2_0_3_reg_1135_pp0_iter47_reg;
            add_i1_2_1_1_reg_1076 <= grp_fu_393_p2;
            add_i1_2_1_2_reg_1141 <= grp_fu_437_p2;
            add_i1_2_1_3_reg_1194 <= grp_fu_473_p2;
            add_i1_2_1_3_reg_1194_pp0_iter49_reg <= add_i1_2_1_3_reg_1194;
            add_i1_2_1_3_reg_1194_pp0_iter50_reg <= add_i1_2_1_3_reg_1194_pp0_iter49_reg;
            add_i1_2_1_3_reg_1194_pp0_iter51_reg <= add_i1_2_1_3_reg_1194_pp0_iter50_reg;
            add_i1_2_1_3_reg_1194_pp0_iter52_reg <= add_i1_2_1_3_reg_1194_pp0_iter51_reg;
            add_i1_2_1_3_reg_1194_pp0_iter53_reg <= add_i1_2_1_3_reg_1194_pp0_iter52_reg;
            add_i1_2_1_3_reg_1194_pp0_iter54_reg <= add_i1_2_1_3_reg_1194_pp0_iter53_reg;
            add_i1_2_1_3_reg_1194_pp0_iter55_reg <= add_i1_2_1_3_reg_1194_pp0_iter54_reg;
            add_i1_2_1_reg_1012 <= grp_fu_360_p2;
            add_i1_2_2_1_reg_1087 <= grp_fu_397_p2;
            add_i1_2_2_2_reg_1146 <= grp_fu_441_p2;
            add_i1_2_2_3_reg_1201 <= grp_fu_477_p2;
            add_i1_2_2_3_reg_1201_pp0_iter49_reg <= add_i1_2_2_3_reg_1201;
            add_i1_2_2_3_reg_1201_pp0_iter50_reg <= add_i1_2_2_3_reg_1201_pp0_iter49_reg;
            add_i1_2_2_3_reg_1201_pp0_iter51_reg <= add_i1_2_2_3_reg_1201_pp0_iter50_reg;
            add_i1_2_2_3_reg_1201_pp0_iter52_reg <= add_i1_2_2_3_reg_1201_pp0_iter51_reg;
            add_i1_2_2_3_reg_1201_pp0_iter53_reg <= add_i1_2_2_3_reg_1201_pp0_iter52_reg;
            add_i1_2_2_3_reg_1201_pp0_iter54_reg <= add_i1_2_2_3_reg_1201_pp0_iter53_reg;
            add_i1_2_2_3_reg_1201_pp0_iter55_reg <= add_i1_2_2_3_reg_1201_pp0_iter54_reg;
            add_i1_2_2_3_reg_1201_pp0_iter56_reg <= add_i1_2_2_3_reg_1201_pp0_iter55_reg;
            add_i1_2_2_3_reg_1201_pp0_iter57_reg <= add_i1_2_2_3_reg_1201_pp0_iter56_reg;
            add_i1_2_2_3_reg_1201_pp0_iter58_reg <= add_i1_2_2_3_reg_1201_pp0_iter57_reg;
            add_i1_2_2_3_reg_1201_pp0_iter59_reg <= add_i1_2_2_3_reg_1201_pp0_iter58_reg;
            add_i1_2_2_3_reg_1201_pp0_iter60_reg <= add_i1_2_2_3_reg_1201_pp0_iter59_reg;
            add_i1_2_2_3_reg_1201_pp0_iter61_reg <= add_i1_2_2_3_reg_1201_pp0_iter60_reg;
            add_i1_2_2_3_reg_1201_pp0_iter62_reg <= add_i1_2_2_3_reg_1201_pp0_iter61_reg;
            add_i1_2_3_2_reg_1151 <= grp_fu_445_p2;
            add_i1_2_3_3_reg_1207 <= grp_fu_481_p2;
            add_i1_2_3_3_reg_1207_pp0_iter49_reg <= add_i1_2_3_3_reg_1207;
            add_i1_2_3_3_reg_1207_pp0_iter50_reg <= add_i1_2_3_3_reg_1207_pp0_iter49_reg;
            add_i1_2_3_3_reg_1207_pp0_iter51_reg <= add_i1_2_3_3_reg_1207_pp0_iter50_reg;
            add_i1_2_3_3_reg_1207_pp0_iter52_reg <= add_i1_2_3_3_reg_1207_pp0_iter51_reg;
            add_i1_2_3_3_reg_1207_pp0_iter53_reg <= add_i1_2_3_3_reg_1207_pp0_iter52_reg;
            add_i1_2_3_3_reg_1207_pp0_iter54_reg <= add_i1_2_3_3_reg_1207_pp0_iter53_reg;
            add_i1_2_3_3_reg_1207_pp0_iter55_reg <= add_i1_2_3_3_reg_1207_pp0_iter54_reg;
            add_i1_2_3_3_reg_1207_pp0_iter56_reg <= add_i1_2_3_3_reg_1207_pp0_iter55_reg;
            add_i1_2_3_3_reg_1207_pp0_iter57_reg <= add_i1_2_3_3_reg_1207_pp0_iter56_reg;
            add_i1_2_3_3_reg_1207_pp0_iter58_reg <= add_i1_2_3_3_reg_1207_pp0_iter57_reg;
            add_i1_2_3_3_reg_1207_pp0_iter59_reg <= add_i1_2_3_3_reg_1207_pp0_iter58_reg;
            add_i1_2_3_3_reg_1207_pp0_iter60_reg <= add_i1_2_3_3_reg_1207_pp0_iter59_reg;
            add_i1_2_3_3_reg_1207_pp0_iter61_reg <= add_i1_2_3_3_reg_1207_pp0_iter60_reg;
            add_i1_2_3_3_reg_1207_pp0_iter62_reg <= add_i1_2_3_3_reg_1207_pp0_iter61_reg;
            add_i1_2_3_3_reg_1207_pp0_iter63_reg <= add_i1_2_3_3_reg_1207_pp0_iter62_reg;
            add_i1_2_3_3_reg_1207_pp0_iter64_reg <= add_i1_2_3_3_reg_1207_pp0_iter63_reg;
            add_i1_2_3_3_reg_1207_pp0_iter65_reg <= add_i1_2_3_3_reg_1207_pp0_iter64_reg;
            add_i1_2_3_3_reg_1207_pp0_iter66_reg <= add_i1_2_3_3_reg_1207_pp0_iter65_reg;
            add_i1_2_3_3_reg_1207_pp0_iter67_reg <= add_i1_2_3_3_reg_1207_pp0_iter66_reg;
            add_i1_2_3_3_reg_1207_pp0_iter68_reg <= add_i1_2_3_3_reg_1207_pp0_iter67_reg;
            add_i1_2_3_3_reg_1207_pp0_iter69_reg <= add_i1_2_3_3_reg_1207_pp0_iter68_reg;
            add_i1_reg_914 <= grp_fu_318_p2;
            add_i2_0_0_1_reg_1297 <= grp_fu_515_p2;
            add_i2_0_0_2_reg_1378 <= grp_fu_563_p2;
            add_i2_0_0_3_reg_1459 <= grp_fu_611_p2;
            add_i2_0_1_1_reg_1309 <= grp_fu_519_p2;
            add_i2_0_1_2_reg_1390 <= grp_fu_567_p2;
            add_i2_0_1_3_reg_1464 <= grp_fu_615_p2;
            add_i2_0_1_reg_1239 <= grp_fu_490_p2;
            add_i2_0_2_1_reg_1314 <= grp_fu_523_p2;
            add_i2_0_2_2_reg_1395 <= grp_fu_571_p2;
            add_i2_0_2_3_reg_1469 <= grp_fu_619_p2;
            add_i2_0_3_1_reg_1319 <= grp_fu_527_p2;
            add_i2_0_3_2_reg_1400 <= grp_fu_575_p2;
            add_i2_0_3_3_reg_1474 <= grp_fu_623_p2;
            add_i2_1_0_1_reg_1324 <= grp_fu_531_p2;
            add_i2_1_0_2_reg_1405 <= grp_fu_579_p2;
            add_i2_1_0_3_reg_1479 <= grp_fu_627_p2;
            add_i2_1_1_1_reg_1336 <= grp_fu_535_p2;
            add_i2_1_1_2_reg_1417 <= grp_fu_583_p2;
            add_i2_1_1_3_reg_1484 <= grp_fu_631_p2;
            add_i2_1_1_reg_1262 <= grp_fu_500_p2;
            add_i2_1_2_1_reg_1341 <= grp_fu_539_p2;
            add_i2_1_2_2_reg_1422 <= grp_fu_587_p2;
            add_i2_1_2_3_reg_1489 <= grp_fu_635_p2;
            add_i2_1_3_1_reg_1346 <= grp_fu_543_p2;
            add_i2_1_3_2_reg_1427 <= grp_fu_591_p2;
            add_i2_1_3_3_reg_1494 <= grp_fu_639_p2;
            add_i2_1_reg_1251 <= grp_fu_495_p2;
            add_i2_2_0_1_reg_1351 <= grp_fu_547_p2;
            add_i2_2_0_2_reg_1432 <= grp_fu_595_p2;
            add_i2_2_0_3_reg_1499 <= grp_fu_643_p2;
            add_i2_2_1_1_reg_1363 <= grp_fu_551_p2;
            add_i2_2_1_2_reg_1444 <= grp_fu_599_p2;
            add_i2_2_1_3_reg_1504 <= grp_fu_647_p2;
            add_i2_2_1_reg_1285 <= grp_fu_510_p2;
            add_i2_2_2_1_reg_1368 <= grp_fu_555_p2;
            add_i2_2_2_2_reg_1449 <= grp_fu_603_p2;
            add_i2_2_2_3_reg_1509 <= grp_fu_651_p2;
            add_i2_2_3_1_reg_1373 <= grp_fu_559_p2;
            add_i2_2_3_2_reg_1454 <= grp_fu_607_p2;
            add_i2_2_3_3_reg_1514 <= grp_fu_655_p2;
            add_i2_2_reg_1274 <= grp_fu_505_p2;
            add_i2_reg_1228 <= grp_fu_485_p2;
            add_i_0_0_3_reg_872 <= grp_fu_288_p2;
            add_i_0_1_3_reg_878 <= grp_fu_293_p2;
            add_i_0_1_3_reg_878_pp0_iter14_reg <= add_i_0_1_3_reg_878;
            add_i_0_1_3_reg_878_pp0_iter15_reg <= add_i_0_1_3_reg_878_pp0_iter14_reg;
            add_i_0_1_3_reg_878_pp0_iter16_reg <= add_i_0_1_3_reg_878_pp0_iter15_reg;
            add_i_0_1_3_reg_878_pp0_iter17_reg <= add_i_0_1_3_reg_878_pp0_iter16_reg;
            add_i_0_1_3_reg_878_pp0_iter18_reg <= add_i_0_1_3_reg_878_pp0_iter17_reg;
            add_i_0_1_3_reg_878_pp0_iter19_reg <= add_i_0_1_3_reg_878_pp0_iter18_reg;
            add_i_0_1_3_reg_878_pp0_iter20_reg <= add_i_0_1_3_reg_878_pp0_iter19_reg;
            add_i_0_1_3_reg_878_pp0_iter21_reg <= add_i_0_1_3_reg_878_pp0_iter20_reg;
            add_i_0_1_3_reg_878_pp0_iter22_reg <= add_i_0_1_3_reg_878_pp0_iter21_reg;
            add_i_0_1_3_reg_878_pp0_iter23_reg <= add_i_0_1_3_reg_878_pp0_iter22_reg;
            add_i_0_1_3_reg_878_pp0_iter24_reg <= add_i_0_1_3_reg_878_pp0_iter23_reg;
            add_i_0_1_3_reg_878_pp0_iter25_reg <= add_i_0_1_3_reg_878_pp0_iter24_reg;
            add_i_0_1_3_reg_878_pp0_iter26_reg <= add_i_0_1_3_reg_878_pp0_iter25_reg;
            add_i_0_1_3_reg_878_pp0_iter27_reg <= add_i_0_1_3_reg_878_pp0_iter26_reg;
            add_i_0_1_3_reg_878_pp0_iter28_reg <= add_i_0_1_3_reg_878_pp0_iter27_reg;
            add_i_0_1_3_reg_878_pp0_iter29_reg <= add_i_0_1_3_reg_878_pp0_iter28_reg;
            add_i_0_1_3_reg_878_pp0_iter30_reg <= add_i_0_1_3_reg_878_pp0_iter29_reg;
            add_i_0_1_3_reg_878_pp0_iter31_reg <= add_i_0_1_3_reg_878_pp0_iter30_reg;
            add_i_0_1_3_reg_878_pp0_iter32_reg <= add_i_0_1_3_reg_878_pp0_iter31_reg;
            add_i_0_1_3_reg_878_pp0_iter33_reg <= add_i_0_1_3_reg_878_pp0_iter32_reg;
            add_i_0_1_3_reg_878_pp0_iter34_reg <= add_i_0_1_3_reg_878_pp0_iter33_reg;
            add_i_0_3_3_reg_952 <= grp_fu_323_p2;
            add_i_0_3_3_reg_952_pp0_iter28_reg <= add_i_0_3_3_reg_952;
            add_i_0_3_3_reg_952_pp0_iter29_reg <= add_i_0_3_3_reg_952_pp0_iter28_reg;
            add_i_0_3_3_reg_952_pp0_iter30_reg <= add_i_0_3_3_reg_952_pp0_iter29_reg;
            add_i_0_3_3_reg_952_pp0_iter31_reg <= add_i_0_3_3_reg_952_pp0_iter30_reg;
            add_i_0_3_3_reg_952_pp0_iter32_reg <= add_i_0_3_3_reg_952_pp0_iter31_reg;
            add_i_0_3_3_reg_952_pp0_iter33_reg <= add_i_0_3_3_reg_952_pp0_iter32_reg;
            add_i_0_3_3_reg_952_pp0_iter34_reg <= add_i_0_3_3_reg_952_pp0_iter33_reg;
            add_i_0_3_3_reg_952_pp0_iter35_reg <= add_i_0_3_3_reg_952_pp0_iter34_reg;
            add_i_0_3_3_reg_952_pp0_iter36_reg <= add_i_0_3_3_reg_952_pp0_iter35_reg;
            add_i_0_3_3_reg_952_pp0_iter37_reg <= add_i_0_3_3_reg_952_pp0_iter36_reg;
            add_i_0_3_3_reg_952_pp0_iter38_reg <= add_i_0_3_3_reg_952_pp0_iter37_reg;
            add_i_0_3_3_reg_952_pp0_iter39_reg <= add_i_0_3_3_reg_952_pp0_iter38_reg;
            add_i_0_3_3_reg_952_pp0_iter40_reg <= add_i_0_3_3_reg_952_pp0_iter39_reg;
            add_i_0_3_3_reg_952_pp0_iter41_reg <= add_i_0_3_3_reg_952_pp0_iter40_reg;
            add_i_1_0_3_reg_886 <= grp_fu_298_p2;
            add_i_1_0_3_reg_886_pp0_iter14_reg <= add_i_1_0_3_reg_886;
            add_i_1_0_3_reg_886_pp0_iter15_reg <= add_i_1_0_3_reg_886_pp0_iter14_reg;
            add_i_1_0_3_reg_886_pp0_iter16_reg <= add_i_1_0_3_reg_886_pp0_iter15_reg;
            add_i_1_0_3_reg_886_pp0_iter17_reg <= add_i_1_0_3_reg_886_pp0_iter16_reg;
            add_i_1_0_3_reg_886_pp0_iter18_reg <= add_i_1_0_3_reg_886_pp0_iter17_reg;
            add_i_1_0_3_reg_886_pp0_iter19_reg <= add_i_1_0_3_reg_886_pp0_iter18_reg;
            add_i_1_0_3_reg_886_pp0_iter20_reg <= add_i_1_0_3_reg_886_pp0_iter19_reg;
            add_i_1_0_3_reg_886_pp0_iter21_reg <= add_i_1_0_3_reg_886_pp0_iter20_reg;
            add_i_1_0_3_reg_886_pp0_iter22_reg <= add_i_1_0_3_reg_886_pp0_iter21_reg;
            add_i_1_0_3_reg_886_pp0_iter23_reg <= add_i_1_0_3_reg_886_pp0_iter22_reg;
            add_i_1_0_3_reg_886_pp0_iter24_reg <= add_i_1_0_3_reg_886_pp0_iter23_reg;
            add_i_1_0_3_reg_886_pp0_iter25_reg <= add_i_1_0_3_reg_886_pp0_iter24_reg;
            add_i_1_0_3_reg_886_pp0_iter26_reg <= add_i_1_0_3_reg_886_pp0_iter25_reg;
            add_i_1_0_3_reg_886_pp0_iter27_reg <= add_i_1_0_3_reg_886_pp0_iter26_reg;
            add_i_1_0_3_reg_886_pp0_iter28_reg <= add_i_1_0_3_reg_886_pp0_iter27_reg;
            add_i_1_0_3_reg_886_pp0_iter29_reg <= add_i_1_0_3_reg_886_pp0_iter28_reg;
            add_i_1_0_3_reg_886_pp0_iter30_reg <= add_i_1_0_3_reg_886_pp0_iter29_reg;
            add_i_1_0_3_reg_886_pp0_iter31_reg <= add_i_1_0_3_reg_886_pp0_iter30_reg;
            add_i_1_0_3_reg_886_pp0_iter32_reg <= add_i_1_0_3_reg_886_pp0_iter31_reg;
            add_i_1_0_3_reg_886_pp0_iter33_reg <= add_i_1_0_3_reg_886_pp0_iter32_reg;
            add_i_1_0_3_reg_886_pp0_iter34_reg <= add_i_1_0_3_reg_886_pp0_iter33_reg;
            add_i_1_1_3_reg_894 <= grp_fu_303_p2;
            add_i_1_1_3_reg_894_pp0_iter14_reg <= add_i_1_1_3_reg_894;
            add_i_1_1_3_reg_894_pp0_iter15_reg <= add_i_1_1_3_reg_894_pp0_iter14_reg;
            add_i_1_1_3_reg_894_pp0_iter16_reg <= add_i_1_1_3_reg_894_pp0_iter15_reg;
            add_i_1_1_3_reg_894_pp0_iter17_reg <= add_i_1_1_3_reg_894_pp0_iter16_reg;
            add_i_1_1_3_reg_894_pp0_iter18_reg <= add_i_1_1_3_reg_894_pp0_iter17_reg;
            add_i_1_1_3_reg_894_pp0_iter19_reg <= add_i_1_1_3_reg_894_pp0_iter18_reg;
            add_i_1_1_3_reg_894_pp0_iter20_reg <= add_i_1_1_3_reg_894_pp0_iter19_reg;
            add_i_1_1_3_reg_894_pp0_iter21_reg <= add_i_1_1_3_reg_894_pp0_iter20_reg;
            add_i_1_1_3_reg_894_pp0_iter22_reg <= add_i_1_1_3_reg_894_pp0_iter21_reg;
            add_i_1_1_3_reg_894_pp0_iter23_reg <= add_i_1_1_3_reg_894_pp0_iter22_reg;
            add_i_1_1_3_reg_894_pp0_iter24_reg <= add_i_1_1_3_reg_894_pp0_iter23_reg;
            add_i_1_1_3_reg_894_pp0_iter25_reg <= add_i_1_1_3_reg_894_pp0_iter24_reg;
            add_i_1_1_3_reg_894_pp0_iter26_reg <= add_i_1_1_3_reg_894_pp0_iter25_reg;
            add_i_1_1_3_reg_894_pp0_iter27_reg <= add_i_1_1_3_reg_894_pp0_iter26_reg;
            add_i_1_3_3_reg_958 <= grp_fu_328_p2;
            add_i_1_3_3_reg_958_pp0_iter28_reg <= add_i_1_3_3_reg_958;
            add_i_1_3_3_reg_958_pp0_iter29_reg <= add_i_1_3_3_reg_958_pp0_iter28_reg;
            add_i_1_3_3_reg_958_pp0_iter30_reg <= add_i_1_3_3_reg_958_pp0_iter29_reg;
            add_i_1_3_3_reg_958_pp0_iter31_reg <= add_i_1_3_3_reg_958_pp0_iter30_reg;
            add_i_1_3_3_reg_958_pp0_iter32_reg <= add_i_1_3_3_reg_958_pp0_iter31_reg;
            add_i_1_3_3_reg_958_pp0_iter33_reg <= add_i_1_3_3_reg_958_pp0_iter32_reg;
            add_i_1_3_3_reg_958_pp0_iter34_reg <= add_i_1_3_3_reg_958_pp0_iter33_reg;
            add_i_1_3_3_reg_958_pp0_iter35_reg <= add_i_1_3_3_reg_958_pp0_iter34_reg;
            add_i_1_3_3_reg_958_pp0_iter36_reg <= add_i_1_3_3_reg_958_pp0_iter35_reg;
            add_i_1_3_3_reg_958_pp0_iter37_reg <= add_i_1_3_3_reg_958_pp0_iter36_reg;
            add_i_1_3_3_reg_958_pp0_iter38_reg <= add_i_1_3_3_reg_958_pp0_iter37_reg;
            add_i_1_3_3_reg_958_pp0_iter39_reg <= add_i_1_3_3_reg_958_pp0_iter38_reg;
            add_i_1_3_3_reg_958_pp0_iter40_reg <= add_i_1_3_3_reg_958_pp0_iter39_reg;
            add_i_1_3_3_reg_958_pp0_iter41_reg <= add_i_1_3_3_reg_958_pp0_iter40_reg;
            add_i_2_0_3_reg_900 <= grp_fu_308_p2;
            add_i_2_0_3_reg_900_pp0_iter14_reg <= add_i_2_0_3_reg_900;
            add_i_2_0_3_reg_900_pp0_iter15_reg <= add_i_2_0_3_reg_900_pp0_iter14_reg;
            add_i_2_0_3_reg_900_pp0_iter16_reg <= add_i_2_0_3_reg_900_pp0_iter15_reg;
            add_i_2_0_3_reg_900_pp0_iter17_reg <= add_i_2_0_3_reg_900_pp0_iter16_reg;
            add_i_2_0_3_reg_900_pp0_iter18_reg <= add_i_2_0_3_reg_900_pp0_iter17_reg;
            add_i_2_0_3_reg_900_pp0_iter19_reg <= add_i_2_0_3_reg_900_pp0_iter18_reg;
            add_i_2_0_3_reg_900_pp0_iter20_reg <= add_i_2_0_3_reg_900_pp0_iter19_reg;
            add_i_2_0_3_reg_900_pp0_iter21_reg <= add_i_2_0_3_reg_900_pp0_iter20_reg;
            add_i_2_0_3_reg_900_pp0_iter22_reg <= add_i_2_0_3_reg_900_pp0_iter21_reg;
            add_i_2_0_3_reg_900_pp0_iter23_reg <= add_i_2_0_3_reg_900_pp0_iter22_reg;
            add_i_2_0_3_reg_900_pp0_iter24_reg <= add_i_2_0_3_reg_900_pp0_iter23_reg;
            add_i_2_0_3_reg_900_pp0_iter25_reg <= add_i_2_0_3_reg_900_pp0_iter24_reg;
            add_i_2_0_3_reg_900_pp0_iter26_reg <= add_i_2_0_3_reg_900_pp0_iter25_reg;
            add_i_2_0_3_reg_900_pp0_iter27_reg <= add_i_2_0_3_reg_900_pp0_iter26_reg;
            add_i_2_2_3_reg_907 <= grp_fu_313_p2;
            add_i_2_2_3_reg_907_pp0_iter21_reg <= add_i_2_2_3_reg_907;
            add_i_2_2_3_reg_907_pp0_iter22_reg <= add_i_2_2_3_reg_907_pp0_iter21_reg;
            add_i_2_2_3_reg_907_pp0_iter23_reg <= add_i_2_2_3_reg_907_pp0_iter22_reg;
            add_i_2_2_3_reg_907_pp0_iter24_reg <= add_i_2_2_3_reg_907_pp0_iter23_reg;
            add_i_2_2_3_reg_907_pp0_iter25_reg <= add_i_2_2_3_reg_907_pp0_iter24_reg;
            add_i_2_2_3_reg_907_pp0_iter26_reg <= add_i_2_2_3_reg_907_pp0_iter25_reg;
            add_i_2_2_3_reg_907_pp0_iter27_reg <= add_i_2_2_3_reg_907_pp0_iter26_reg;
            add_i_2_2_3_reg_907_pp0_iter28_reg <= add_i_2_2_3_reg_907_pp0_iter27_reg;
            add_i_2_2_3_reg_907_pp0_iter29_reg <= add_i_2_2_3_reg_907_pp0_iter28_reg;
            add_i_2_2_3_reg_907_pp0_iter30_reg <= add_i_2_2_3_reg_907_pp0_iter29_reg;
            add_i_2_2_3_reg_907_pp0_iter31_reg <= add_i_2_2_3_reg_907_pp0_iter30_reg;
            add_i_2_2_3_reg_907_pp0_iter32_reg <= add_i_2_2_3_reg_907_pp0_iter31_reg;
            add_i_2_2_3_reg_907_pp0_iter33_reg <= add_i_2_2_3_reg_907_pp0_iter32_reg;
            add_i_2_2_3_reg_907_pp0_iter34_reg <= add_i_2_2_3_reg_907_pp0_iter33_reg;
            add_i_2_3_3_reg_964 <= grp_fu_333_p2;
            add_i_2_3_3_reg_964_pp0_iter28_reg <= add_i_2_3_3_reg_964;
            add_i_2_3_3_reg_964_pp0_iter29_reg <= add_i_2_3_3_reg_964_pp0_iter28_reg;
            add_i_2_3_3_reg_964_pp0_iter30_reg <= add_i_2_3_3_reg_964_pp0_iter29_reg;
            add_i_2_3_3_reg_964_pp0_iter31_reg <= add_i_2_3_3_reg_964_pp0_iter30_reg;
            add_i_2_3_3_reg_964_pp0_iter32_reg <= add_i_2_3_3_reg_964_pp0_iter31_reg;
            add_i_2_3_3_reg_964_pp0_iter33_reg <= add_i_2_3_3_reg_964_pp0_iter32_reg;
            add_i_2_3_3_reg_964_pp0_iter34_reg <= add_i_2_3_3_reg_964_pp0_iter33_reg;
            add_i_2_3_3_reg_964_pp0_iter35_reg <= add_i_2_3_3_reg_964_pp0_iter34_reg;
            add_i_2_3_3_reg_964_pp0_iter36_reg <= add_i_2_3_3_reg_964_pp0_iter35_reg;
            add_i_2_3_3_reg_964_pp0_iter37_reg <= add_i_2_3_3_reg_964_pp0_iter36_reg;
            add_i_2_3_3_reg_964_pp0_iter38_reg <= add_i_2_3_3_reg_964_pp0_iter37_reg;
            add_i_2_3_3_reg_964_pp0_iter39_reg <= add_i_2_3_3_reg_964_pp0_iter38_reg;
            add_i_2_3_3_reg_964_pp0_iter40_reg <= add_i_2_3_3_reg_964_pp0_iter39_reg;
            add_i_2_3_3_reg_964_pp0_iter41_reg <= add_i_2_3_3_reg_964_pp0_iter40_reg;
            mul_i1_0_0_1_reg_919 <= grp_fu_677_p2;
            mul_i1_0_0_1_reg_919_pp0_iter21_reg <= mul_i1_0_0_1_reg_919;
            mul_i1_0_0_1_reg_919_pp0_iter22_reg <= mul_i1_0_0_1_reg_919_pp0_iter21_reg;
            mul_i1_0_0_1_reg_919_pp0_iter23_reg <= mul_i1_0_0_1_reg_919_pp0_iter22_reg;
            mul_i1_0_0_1_reg_919_pp0_iter24_reg <= mul_i1_0_0_1_reg_919_pp0_iter23_reg;
            mul_i1_0_0_1_reg_919_pp0_iter25_reg <= mul_i1_0_0_1_reg_919_pp0_iter24_reg;
            mul_i1_0_0_1_reg_919_pp0_iter26_reg <= mul_i1_0_0_1_reg_919_pp0_iter25_reg;
            mul_i1_0_0_1_reg_919_pp0_iter27_reg <= mul_i1_0_0_1_reg_919_pp0_iter26_reg;
            mul_i1_0_0_1_reg_919_pp0_iter28_reg <= mul_i1_0_0_1_reg_919_pp0_iter27_reg;
            mul_i1_0_0_1_reg_919_pp0_iter29_reg <= mul_i1_0_0_1_reg_919_pp0_iter28_reg;
            mul_i1_0_0_1_reg_919_pp0_iter30_reg <= mul_i1_0_0_1_reg_919_pp0_iter29_reg;
            mul_i1_0_0_1_reg_919_pp0_iter31_reg <= mul_i1_0_0_1_reg_919_pp0_iter30_reg;
            mul_i1_0_0_1_reg_919_pp0_iter32_reg <= mul_i1_0_0_1_reg_919_pp0_iter31_reg;
            mul_i1_0_0_1_reg_919_pp0_iter33_reg <= mul_i1_0_0_1_reg_919_pp0_iter32_reg;
            mul_i1_0_0_1_reg_919_pp0_iter34_reg <= mul_i1_0_0_1_reg_919_pp0_iter33_reg;
            mul_i1_0_0_2_reg_975 <= grp_fu_702_p2;
            mul_i1_0_0_3_reg_1023 <= grp_fu_717_p2;
            mul_i1_0_0_3_reg_1023_pp0_iter35_reg <= mul_i1_0_0_3_reg_1023;
            mul_i1_0_0_3_reg_1023_pp0_iter36_reg <= mul_i1_0_0_3_reg_1023_pp0_iter35_reg;
            mul_i1_0_0_3_reg_1023_pp0_iter37_reg <= mul_i1_0_0_3_reg_1023_pp0_iter36_reg;
            mul_i1_0_0_3_reg_1023_pp0_iter38_reg <= mul_i1_0_0_3_reg_1023_pp0_iter37_reg;
            mul_i1_0_0_3_reg_1023_pp0_iter39_reg <= mul_i1_0_0_3_reg_1023_pp0_iter38_reg;
            mul_i1_0_0_3_reg_1023_pp0_iter40_reg <= mul_i1_0_0_3_reg_1023_pp0_iter39_reg;
            mul_i1_0_0_3_reg_1023_pp0_iter41_reg <= mul_i1_0_0_3_reg_1023_pp0_iter40_reg;
            mul_i1_0_1_reg_927 <= grp_fu_682_p2;
            mul_i1_1_0_1_reg_932 <= grp_fu_687_p2;
            mul_i1_1_0_1_reg_932_pp0_iter21_reg <= mul_i1_1_0_1_reg_932;
            mul_i1_1_0_1_reg_932_pp0_iter22_reg <= mul_i1_1_0_1_reg_932_pp0_iter21_reg;
            mul_i1_1_0_1_reg_932_pp0_iter23_reg <= mul_i1_1_0_1_reg_932_pp0_iter22_reg;
            mul_i1_1_0_1_reg_932_pp0_iter24_reg <= mul_i1_1_0_1_reg_932_pp0_iter23_reg;
            mul_i1_1_0_1_reg_932_pp0_iter25_reg <= mul_i1_1_0_1_reg_932_pp0_iter24_reg;
            mul_i1_1_0_1_reg_932_pp0_iter26_reg <= mul_i1_1_0_1_reg_932_pp0_iter25_reg;
            mul_i1_1_0_1_reg_932_pp0_iter27_reg <= mul_i1_1_0_1_reg_932_pp0_iter26_reg;
            mul_i1_1_0_2_reg_991 <= grp_fu_707_p2;
            mul_i1_1_0_3_reg_1046 <= grp_fu_722_p2;
            mul_i1_1_0_3_reg_1046_pp0_iter35_reg <= mul_i1_1_0_3_reg_1046;
            mul_i1_1_0_3_reg_1046_pp0_iter36_reg <= mul_i1_1_0_3_reg_1046_pp0_iter35_reg;
            mul_i1_1_0_3_reg_1046_pp0_iter37_reg <= mul_i1_1_0_3_reg_1046_pp0_iter36_reg;
            mul_i1_1_0_3_reg_1046_pp0_iter38_reg <= mul_i1_1_0_3_reg_1046_pp0_iter37_reg;
            mul_i1_1_0_3_reg_1046_pp0_iter39_reg <= mul_i1_1_0_3_reg_1046_pp0_iter38_reg;
            mul_i1_1_0_3_reg_1046_pp0_iter40_reg <= mul_i1_1_0_3_reg_1046_pp0_iter39_reg;
            mul_i1_1_0_3_reg_1046_pp0_iter41_reg <= mul_i1_1_0_3_reg_1046_pp0_iter40_reg;
            mul_i1_1_1_reg_938 <= grp_fu_692_p2;
            mul_i1_1_1_reg_938_pp0_iter21_reg <= mul_i1_1_1_reg_938;
            mul_i1_1_1_reg_938_pp0_iter22_reg <= mul_i1_1_1_reg_938_pp0_iter21_reg;
            mul_i1_1_1_reg_938_pp0_iter23_reg <= mul_i1_1_1_reg_938_pp0_iter22_reg;
            mul_i1_1_1_reg_938_pp0_iter24_reg <= mul_i1_1_1_reg_938_pp0_iter23_reg;
            mul_i1_1_1_reg_938_pp0_iter25_reg <= mul_i1_1_1_reg_938_pp0_iter24_reg;
            mul_i1_1_1_reg_938_pp0_iter26_reg <= mul_i1_1_1_reg_938_pp0_iter25_reg;
            mul_i1_1_1_reg_938_pp0_iter27_reg <= mul_i1_1_1_reg_938_pp0_iter26_reg;
            mul_i1_1_1_reg_938_pp0_iter28_reg <= mul_i1_1_1_reg_938_pp0_iter27_reg;
            mul_i1_1_1_reg_938_pp0_iter29_reg <= mul_i1_1_1_reg_938_pp0_iter28_reg;
            mul_i1_1_1_reg_938_pp0_iter30_reg <= mul_i1_1_1_reg_938_pp0_iter29_reg;
            mul_i1_1_1_reg_938_pp0_iter31_reg <= mul_i1_1_1_reg_938_pp0_iter30_reg;
            mul_i1_1_1_reg_938_pp0_iter32_reg <= mul_i1_1_1_reg_938_pp0_iter31_reg;
            mul_i1_1_1_reg_938_pp0_iter33_reg <= mul_i1_1_1_reg_938_pp0_iter32_reg;
            mul_i1_1_1_reg_938_pp0_iter34_reg <= mul_i1_1_1_reg_938_pp0_iter33_reg;
            mul_i1_2_0_1_reg_945 <= grp_fu_697_p2;
            mul_i1_2_0_1_reg_945_pp0_iter21_reg <= mul_i1_2_0_1_reg_945;
            mul_i1_2_0_1_reg_945_pp0_iter22_reg <= mul_i1_2_0_1_reg_945_pp0_iter21_reg;
            mul_i1_2_0_1_reg_945_pp0_iter23_reg <= mul_i1_2_0_1_reg_945_pp0_iter22_reg;
            mul_i1_2_0_1_reg_945_pp0_iter24_reg <= mul_i1_2_0_1_reg_945_pp0_iter23_reg;
            mul_i1_2_0_1_reg_945_pp0_iter25_reg <= mul_i1_2_0_1_reg_945_pp0_iter24_reg;
            mul_i1_2_0_1_reg_945_pp0_iter26_reg <= mul_i1_2_0_1_reg_945_pp0_iter25_reg;
            mul_i1_2_0_1_reg_945_pp0_iter27_reg <= mul_i1_2_0_1_reg_945_pp0_iter26_reg;
            mul_i1_2_0_2_reg_1007 <= grp_fu_712_p2;
            mul_i1_2_0_3_reg_1069 <= grp_fu_727_p2;
            mul_i1_2_0_3_reg_1069_pp0_iter35_reg <= mul_i1_2_0_3_reg_1069;
            mul_i1_2_0_3_reg_1069_pp0_iter36_reg <= mul_i1_2_0_3_reg_1069_pp0_iter35_reg;
            mul_i1_2_0_3_reg_1069_pp0_iter37_reg <= mul_i1_2_0_3_reg_1069_pp0_iter36_reg;
            mul_i1_2_0_3_reg_1069_pp0_iter38_reg <= mul_i1_2_0_3_reg_1069_pp0_iter37_reg;
            mul_i1_2_0_3_reg_1069_pp0_iter39_reg <= mul_i1_2_0_3_reg_1069_pp0_iter38_reg;
            mul_i1_2_0_3_reg_1069_pp0_iter40_reg <= mul_i1_2_0_3_reg_1069_pp0_iter39_reg;
            mul_i1_2_0_3_reg_1069_pp0_iter41_reg <= mul_i1_2_0_3_reg_1069_pp0_iter40_reg;
            mul_i1_2_1_2_reg_1081 <= grp_fu_732_p2;
            mul_i2_0_0_1_reg_1233 <= grp_fu_752_p2;
            mul_i2_0_0_2_reg_1302 <= grp_fu_782_p2;
            mul_i2_0_0_3_reg_1383 <= grp_fu_797_p2;
            mul_i2_0_1_reg_1213 <= grp_fu_737_p2;
            mul_i2_0_2_1_reg_1246 <= grp_fu_757_p2;
            mul_i2_1_0_1_reg_1256 <= grp_fu_762_p2;
            mul_i2_1_0_2_reg_1329 <= grp_fu_787_p2;
            mul_i2_1_0_3_reg_1410 <= grp_fu_802_p2;
            mul_i2_1_1_reg_1218 <= grp_fu_742_p2;
            mul_i2_1_2_1_reg_1269 <= grp_fu_767_p2;
            mul_i2_2_0_1_reg_1279 <= grp_fu_772_p2;
            mul_i2_2_0_2_reg_1356 <= grp_fu_792_p2;
            mul_i2_2_0_3_reg_1437 <= grp_fu_807_p2;
            mul_i2_2_1_reg_1223 <= grp_fu_747_p2;
            mul_i2_2_2_1_reg_1292 <= grp_fu_777_p2;
            mul_i_0_0_3_reg_854 <= grp_fu_659_p2;
            mul_i_1_0_3_reg_860 <= grp_fu_665_p2;
            mul_i_2_0_3_reg_866 <= grp_fu_671_p2;
            mul_i_2_0_3_reg_866_pp0_iter10_reg <= mul_i_2_0_3_reg_866_pp0_iter9_reg;
            mul_i_2_0_3_reg_866_pp0_iter11_reg <= mul_i_2_0_3_reg_866_pp0_iter10_reg;
            mul_i_2_0_3_reg_866_pp0_iter12_reg <= mul_i_2_0_3_reg_866_pp0_iter11_reg;
            mul_i_2_0_3_reg_866_pp0_iter13_reg <= mul_i_2_0_3_reg_866_pp0_iter12_reg;
            mul_i_2_0_3_reg_866_pp0_iter7_reg <= mul_i_2_0_3_reg_866;
            mul_i_2_0_3_reg_866_pp0_iter8_reg <= mul_i_2_0_3_reg_866_pp0_iter7_reg;
            mul_i_2_0_3_reg_866_pp0_iter9_reg <= mul_i_2_0_3_reg_866_pp0_iter8_reg;
            x_read_reg_832_pp0_iter10_reg <= x_read_reg_832_pp0_iter9_reg;
            x_read_reg_832_pp0_iter11_reg <= x_read_reg_832_pp0_iter10_reg;
            x_read_reg_832_pp0_iter12_reg <= x_read_reg_832_pp0_iter11_reg;
            x_read_reg_832_pp0_iter13_reg <= x_read_reg_832_pp0_iter12_reg;
            x_read_reg_832_pp0_iter14_reg <= x_read_reg_832_pp0_iter13_reg;
            x_read_reg_832_pp0_iter15_reg <= x_read_reg_832_pp0_iter14_reg;
            x_read_reg_832_pp0_iter16_reg <= x_read_reg_832_pp0_iter15_reg;
            x_read_reg_832_pp0_iter17_reg <= x_read_reg_832_pp0_iter16_reg;
            x_read_reg_832_pp0_iter18_reg <= x_read_reg_832_pp0_iter17_reg;
            x_read_reg_832_pp0_iter19_reg <= x_read_reg_832_pp0_iter18_reg;
            x_read_reg_832_pp0_iter20_reg <= x_read_reg_832_pp0_iter19_reg;
            x_read_reg_832_pp0_iter2_reg <= x_read_reg_832_pp0_iter1_reg;
            x_read_reg_832_pp0_iter3_reg <= x_read_reg_832_pp0_iter2_reg;
            x_read_reg_832_pp0_iter4_reg <= x_read_reg_832_pp0_iter3_reg;
            x_read_reg_832_pp0_iter5_reg <= x_read_reg_832_pp0_iter4_reg;
            x_read_reg_832_pp0_iter6_reg <= x_read_reg_832_pp0_iter5_reg;
            x_read_reg_832_pp0_iter7_reg <= x_read_reg_832_pp0_iter6_reg;
            x_read_reg_832_pp0_iter8_reg <= x_read_reg_832_pp0_iter7_reg;
            x_read_reg_832_pp0_iter9_reg <= x_read_reg_832_pp0_iter8_reg;
            y_read_reg_826_pp0_iter10_reg <= y_read_reg_826_pp0_iter9_reg;
            y_read_reg_826_pp0_iter11_reg <= y_read_reg_826_pp0_iter10_reg;
            y_read_reg_826_pp0_iter12_reg <= y_read_reg_826_pp0_iter11_reg;
            y_read_reg_826_pp0_iter13_reg <= y_read_reg_826_pp0_iter12_reg;
            y_read_reg_826_pp0_iter14_reg <= y_read_reg_826_pp0_iter13_reg;
            y_read_reg_826_pp0_iter15_reg <= y_read_reg_826_pp0_iter14_reg;
            y_read_reg_826_pp0_iter16_reg <= y_read_reg_826_pp0_iter15_reg;
            y_read_reg_826_pp0_iter17_reg <= y_read_reg_826_pp0_iter16_reg;
            y_read_reg_826_pp0_iter18_reg <= y_read_reg_826_pp0_iter17_reg;
            y_read_reg_826_pp0_iter19_reg <= y_read_reg_826_pp0_iter18_reg;
            y_read_reg_826_pp0_iter20_reg <= y_read_reg_826_pp0_iter19_reg;
            y_read_reg_826_pp0_iter2_reg <= y_read_reg_826_pp0_iter1_reg;
            y_read_reg_826_pp0_iter3_reg <= y_read_reg_826_pp0_iter2_reg;
            y_read_reg_826_pp0_iter4_reg <= y_read_reg_826_pp0_iter3_reg;
            y_read_reg_826_pp0_iter5_reg <= y_read_reg_826_pp0_iter4_reg;
            y_read_reg_826_pp0_iter6_reg <= y_read_reg_826_pp0_iter5_reg;
            y_read_reg_826_pp0_iter7_reg <= y_read_reg_826_pp0_iter6_reg;
            y_read_reg_826_pp0_iter8_reg <= y_read_reg_826_pp0_iter7_reg;
            y_read_reg_826_pp0_iter9_reg <= y_read_reg_826_pp0_iter8_reg;
            z_read_reg_820_pp0_iter10_reg <= z_read_reg_820_pp0_iter9_reg;
            z_read_reg_820_pp0_iter11_reg <= z_read_reg_820_pp0_iter10_reg;
            z_read_reg_820_pp0_iter12_reg <= z_read_reg_820_pp0_iter11_reg;
            z_read_reg_820_pp0_iter13_reg <= z_read_reg_820_pp0_iter12_reg;
            z_read_reg_820_pp0_iter14_reg <= z_read_reg_820_pp0_iter13_reg;
            z_read_reg_820_pp0_iter15_reg <= z_read_reg_820_pp0_iter14_reg;
            z_read_reg_820_pp0_iter16_reg <= z_read_reg_820_pp0_iter15_reg;
            z_read_reg_820_pp0_iter17_reg <= z_read_reg_820_pp0_iter16_reg;
            z_read_reg_820_pp0_iter18_reg <= z_read_reg_820_pp0_iter17_reg;
            z_read_reg_820_pp0_iter19_reg <= z_read_reg_820_pp0_iter18_reg;
            z_read_reg_820_pp0_iter20_reg <= z_read_reg_820_pp0_iter19_reg;
            z_read_reg_820_pp0_iter2_reg <= z_read_reg_820_pp0_iter1_reg;
            z_read_reg_820_pp0_iter3_reg <= z_read_reg_820_pp0_iter2_reg;
            z_read_reg_820_pp0_iter4_reg <= z_read_reg_820_pp0_iter3_reg;
            z_read_reg_820_pp0_iter5_reg <= z_read_reg_820_pp0_iter4_reg;
            z_read_reg_820_pp0_iter6_reg <= z_read_reg_820_pp0_iter5_reg;
            z_read_reg_820_pp0_iter7_reg <= z_read_reg_820_pp0_iter6_reg;
            z_read_reg_820_pp0_iter8_reg <= z_read_reg_820_pp0_iter7_reg;
            z_read_reg_820_pp0_iter9_reg <= z_read_reg_820_pp0_iter8_reg;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_0_ce0 = 1'b1;
        end else begin
            H_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_0_we0 = 1'b1;
        end else begin
            H_0_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_1_ce0 = 1'b1;
        end else begin
            H_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_1_we0 = 1'b1;
        end else begin
            H_0_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_2_ce0 = 1'b1;
        end else begin
            H_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_2_we0 = 1'b1;
        end else begin
            H_0_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_3_ce0 = 1'b1;
        end else begin
            H_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_0_3_we0 = 1'b1;
        end else begin
            H_0_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_0_ce0 = 1'b1;
        end else begin
            H_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_0_we0 = 1'b1;
        end else begin
            H_1_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_1_ce0 = 1'b1;
        end else begin
            H_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_1_we0 = 1'b1;
        end else begin
            H_1_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_2_ce0 = 1'b1;
        end else begin
            H_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_2_we0 = 1'b1;
        end else begin
            H_1_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_3_ce0 = 1'b1;
        end else begin
            H_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_1_3_we0 = 1'b1;
        end else begin
            H_1_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_0_ce0 = 1'b1;
        end else begin
            H_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_0_we0 = 1'b1;
        end else begin
            H_2_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_1_ce0 = 1'b1;
        end else begin
            H_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_1_we0 = 1'b1;
        end else begin
            H_2_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_2_ce0 = 1'b1;
        end else begin
            H_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_2_we0 = 1'b1;
        end else begin
            H_2_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_3_ce0 = 1'b1;
        end else begin
            H_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            H_2_3_we0 = 1'b1;
        end else begin
            H_2_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_0_ce0 = 1'b1;
        end else begin
            H_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_0_we0 = 1'b1;
        end else begin
            H_3_0_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_1_ce0 = 1'b1;
        end else begin
            H_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_1_we0 = 1'b1;
        end else begin
            H_3_1_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_2_ce0 = 1'b1;
        end else begin
            H_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_2_we0 = 1'b1;
        end else begin
            H_3_2_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_3_ce0 = 1'b1;
        end else begin
            H_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_3_3_we0 = 1'b1;
        end else begin
            H_3_3_we0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter77 == 1'b1))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter77 == 1'b0) & (ap_enable_reg_pp0_iter76 == 1'b0) & (ap_enable_reg_pp0_iter75 == 1'b0) 
    & (ap_enable_reg_pp0_iter74 == 1'b0) & (ap_enable_reg_pp0_iter73 == 1'b0) & (ap_enable_reg_pp0_iter72 == 1'b0) & (ap_enable_reg_pp0_iter71 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter70 == 1'b0) & (ap_enable_reg_pp0_iter69 == 1'b0) & (ap_enable_reg_pp0_iter68 == 1'b0) & (ap_enable_reg_pp0_iter67 == 1'b0) & (ap_enable_reg_pp0_iter66 == 1'b0) & (ap_enable_reg_pp0_iter65 == 1'b0) & (ap_enable_reg_pp0_iter64 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter63 == 1'b0) & (ap_enable_reg_pp0_iter62 == 1'b0) & (ap_enable_reg_pp0_iter61 == 1'b0) & (ap_enable_reg_pp0_iter60 == 1'b0) & (ap_enable_reg_pp0_iter59 == 1'b0) & (ap_enable_reg_pp0_iter58 == 1'b0) & (ap_enable_reg_pp0_iter57 == 1'b0) & (ap_enable_reg_pp0_iter56 == 1'b0) & (ap_enable_reg_pp0_iter55 == 1'b0) & (ap_enable_reg_pp0_iter54 == 1'b0) & (ap_enable_reg_pp0_iter53 == 1'b0) & (ap_enable_reg_pp0_iter52 == 1'b0) & (ap_enable_reg_pp0_iter51 == 1'b0) & (ap_enable_reg_pp0_iter50 == 1'b0) & (ap_enable_reg_pp0_iter49 
    == 1'b0) & (ap_enable_reg_pp0_iter48 == 1'b0) & (ap_enable_reg_pp0_iter47 == 1'b0) & (ap_enable_reg_pp0_iter46 == 1'b0) & (ap_enable_reg_pp0_iter45 == 1'b0) & (ap_enable_reg_pp0_iter44 == 1'b0) & (ap_enable_reg_pp0_iter43 == 1'b0) & (ap_enable_reg_pp0_iter42 == 1'b0) & (ap_enable_reg_pp0_iter41 == 1'b0) & (ap_enable_reg_pp0_iter40 == 1'b0) & (ap_enable_reg_pp0_iter39 == 1'b0) & (ap_enable_reg_pp0_iter38 == 1'b0) & (ap_enable_reg_pp0_iter37 == 1'b0) & (ap_enable_reg_pp0_iter36 == 1'b0) & (ap_enable_reg_pp0_iter35 == 1'b0) & (ap_enable_reg_pp0_iter34 == 1'b0) & (ap_enable_reg_pp0_iter33 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter76 == 1'b0) & (ap_enable_reg_pp0_iter75 == 1'b0) & (ap_enable_reg_pp0_iter74 == 1'b0) 
    & (ap_enable_reg_pp0_iter73 == 1'b0) & (ap_enable_reg_pp0_iter72 == 1'b0) & (ap_enable_reg_pp0_iter71 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter70 == 1'b0) & (ap_enable_reg_pp0_iter69 == 1'b0) & (ap_enable_reg_pp0_iter68 == 1'b0) & (ap_enable_reg_pp0_iter67 == 1'b0) & (ap_enable_reg_pp0_iter66 == 1'b0) & (ap_enable_reg_pp0_iter65 == 1'b0) & (ap_enable_reg_pp0_iter64 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter63 == 1'b0) & (ap_enable_reg_pp0_iter62 == 1'b0) & (ap_enable_reg_pp0_iter61 == 1'b0) & (ap_enable_reg_pp0_iter60 == 1'b0) & (ap_enable_reg_pp0_iter59 == 1'b0) & (ap_enable_reg_pp0_iter58 == 1'b0) & (ap_enable_reg_pp0_iter57 == 1'b0) & (ap_enable_reg_pp0_iter56 == 1'b0) & (ap_enable_reg_pp0_iter55 == 1'b0) & (ap_enable_reg_pp0_iter54 == 1'b0) & (ap_enable_reg_pp0_iter53 == 1'b0) & (ap_enable_reg_pp0_iter52 == 1'b0) & (ap_enable_reg_pp0_iter51 == 1'b0) & (ap_enable_reg_pp0_iter50 == 1'b0) & (ap_enable_reg_pp0_iter49 == 1'b0) & (ap_enable_reg_pp0_iter48 
    == 1'b0) & (ap_enable_reg_pp0_iter47 == 1'b0) & (ap_enable_reg_pp0_iter46 == 1'b0) & (ap_enable_reg_pp0_iter45 == 1'b0) & (ap_enable_reg_pp0_iter44 == 1'b0) & (ap_enable_reg_pp0_iter43 == 1'b0) & (ap_enable_reg_pp0_iter42 == 1'b0) & (ap_enable_reg_pp0_iter41 == 1'b0) & (ap_enable_reg_pp0_iter40 == 1'b0) & (ap_enable_reg_pp0_iter39 == 1'b0) & (ap_enable_reg_pp0_iter38 == 1'b0) & (ap_enable_reg_pp0_iter37 == 1'b0) & (ap_enable_reg_pp0_iter36 == 1'b0) & (ap_enable_reg_pp0_iter35 == 1'b0) & (ap_enable_reg_pp0_iter34 == 1'b0) & (ap_enable_reg_pp0_iter33 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0_0to76 = 1'b1;
        end else begin
            ap_idle_pp0_0to76 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (ap_idle_pp0_0to76 == 1'b1))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign H_0_0_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_0_0_d0 = add_i2_0_0_3_reg_1459;

    assign H_0_1_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_0_1_d0 = add_i2_0_1_3_reg_1464;

    assign H_0_2_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_0_2_d0 = add_i2_0_2_3_reg_1469;

    assign H_0_3_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_0_3_d0 = add_i2_0_3_3_reg_1474;

    assign H_1_0_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_1_0_d0 = add_i2_1_0_3_reg_1479;

    assign H_1_1_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_1_1_d0 = add_i2_1_1_3_reg_1484;

    assign H_1_2_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_1_2_d0 = add_i2_1_2_3_reg_1489;

    assign H_1_3_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_1_3_d0 = add_i2_1_3_3_reg_1494;

    assign H_2_0_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_2_0_d0 = add_i2_2_0_3_reg_1499;

    assign H_2_1_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_2_1_d0 = add_i2_2_1_3_reg_1504;

    assign H_2_2_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_2_2_d0 = add_i2_2_2_3_reg_1509;

    assign H_2_3_address0 = H_offset_cast_reg_838_pp0_iter76_reg;

    assign H_2_3_d0 = add_i2_2_3_3_reg_1514;

    assign H_3_0_address0 = H_offset_cast_fu_812_p1;

    assign H_3_0_d0 = 64'd0;

    assign H_3_1_address0 = H_offset_cast_fu_812_p1;

    assign H_3_1_d0 = 64'd0;

    assign H_3_2_address0 = H_offset_cast_fu_812_p1;

    assign H_3_2_d0 = 64'd0;

    assign H_3_3_address0 = H_offset_cast_fu_812_p1;

    assign H_3_3_d0 = 64'd4607182418800017408;

    assign H_offset_cast_fu_812_p1 = H_offset;

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start;

    always @(posedge ap_clk) begin
        H_offset_cast_reg_838[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter1_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter2_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter3_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter4_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter5_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter6_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter7_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter8_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter9_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter10_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter11_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter12_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter13_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter14_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter15_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter16_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter17_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter18_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter19_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter20_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter21_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter22_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter23_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter24_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter25_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter26_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter27_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter28_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter29_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter30_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter31_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter32_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter33_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter34_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter35_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter36_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter37_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter38_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter39_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter40_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter41_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter42_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter43_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter44_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter45_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter46_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter47_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter48_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter49_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter50_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter51_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter52_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter53_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter54_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter55_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter56_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter57_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter58_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter59_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter60_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter61_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter62_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter63_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter64_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter65_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter66_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter67_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter68_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter69_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter70_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter71_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter72_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter73_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter74_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter75_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
        H_offset_cast_reg_838_pp0_iter76_reg[63:3] <= 61'b0000000000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_rpyxyzToH_double_1
