/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_main_Pipeline_VITIS_LOOP_69_4 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    l_TBlock_3_3_3_0194_out,
    l_TBlock_3_3_3_0194_out_ap_vld,
    l_TBlock_3_3_2_0193_out,
    l_TBlock_3_3_2_0193_out_ap_vld,
    l_TBlock_3_3_1_0192_out,
    l_TBlock_3_3_1_0192_out_ap_vld,
    l_TBlock_3_3_0_0191_out,
    l_TBlock_3_3_0_0191_out_ap_vld,
    l_TBlock_3_2_3_0190_out,
    l_TBlock_3_2_3_0190_out_ap_vld,
    l_TBlock_3_2_2_0189_out,
    l_TBlock_3_2_2_0189_out_ap_vld,
    l_TBlock_3_2_1_0188_out,
    l_TBlock_3_2_1_0188_out_ap_vld,
    l_TBlock_3_2_0_0187_out,
    l_TBlock_3_2_0_0187_out_ap_vld,
    l_TBlock_3_1_3_0186_out,
    l_TBlock_3_1_3_0186_out_ap_vld,
    l_TBlock_3_1_2_0185_out,
    l_TBlock_3_1_2_0185_out_ap_vld,
    l_TBlock_3_1_1_0184_out,
    l_TBlock_3_1_1_0184_out_ap_vld,
    l_TBlock_3_1_0_0183_out,
    l_TBlock_3_1_0_0183_out_ap_vld,
    l_TBlock_3_0_3_0182_out,
    l_TBlock_3_0_3_0182_out_ap_vld,
    l_TBlock_3_0_2_0181_out,
    l_TBlock_3_0_2_0181_out_ap_vld,
    l_TBlock_3_0_1_0180_out,
    l_TBlock_3_0_1_0180_out_ap_vld,
    l_TBlock_3_0_0_0179_out,
    l_TBlock_3_0_0_0179_out_ap_vld,
    l_TBlock_2_3_3_0178_out,
    l_TBlock_2_3_3_0178_out_ap_vld,
    l_TBlock_2_3_2_0177_out,
    l_TBlock_2_3_2_0177_out_ap_vld,
    l_TBlock_2_3_1_0176_out,
    l_TBlock_2_3_1_0176_out_ap_vld,
    l_TBlock_2_3_0_0175_out,
    l_TBlock_2_3_0_0175_out_ap_vld,
    l_TBlock_2_2_3_0174_out,
    l_TBlock_2_2_3_0174_out_ap_vld,
    l_TBlock_2_2_2_0173_out,
    l_TBlock_2_2_2_0173_out_ap_vld,
    l_TBlock_2_2_1_0172_out,
    l_TBlock_2_2_1_0172_out_ap_vld,
    l_TBlock_2_2_0_0171_out,
    l_TBlock_2_2_0_0171_out_ap_vld,
    l_TBlock_2_1_3_0170_out,
    l_TBlock_2_1_3_0170_out_ap_vld,
    l_TBlock_2_1_2_0169_out,
    l_TBlock_2_1_2_0169_out_ap_vld,
    l_TBlock_2_1_1_0168_out,
    l_TBlock_2_1_1_0168_out_ap_vld,
    l_TBlock_2_1_0_0167_out,
    l_TBlock_2_1_0_0167_out_ap_vld,
    l_TBlock_2_0_3_0166_out,
    l_TBlock_2_0_3_0166_out_ap_vld,
    l_TBlock_2_0_2_0165_out,
    l_TBlock_2_0_2_0165_out_ap_vld,
    l_TBlock_2_0_1_0164_out,
    l_TBlock_2_0_1_0164_out_ap_vld,
    l_TBlock_2_0_0_0163_out,
    l_TBlock_2_0_0_0163_out_ap_vld,
    l_TBlock_1_3_3_0162_out,
    l_TBlock_1_3_3_0162_out_ap_vld,
    l_TBlock_1_3_2_0161_out,
    l_TBlock_1_3_2_0161_out_ap_vld,
    l_TBlock_1_3_1_0160_out,
    l_TBlock_1_3_1_0160_out_ap_vld,
    l_TBlock_1_3_0_0159_out,
    l_TBlock_1_3_0_0159_out_ap_vld,
    l_TBlock_1_2_3_0158_out,
    l_TBlock_1_2_3_0158_out_ap_vld,
    l_TBlock_1_2_2_0157_out,
    l_TBlock_1_2_2_0157_out_ap_vld,
    l_TBlock_1_2_1_0156_out,
    l_TBlock_1_2_1_0156_out_ap_vld,
    l_TBlock_1_2_0_0155_out,
    l_TBlock_1_2_0_0155_out_ap_vld,
    l_TBlock_1_1_3_0154_out,
    l_TBlock_1_1_3_0154_out_ap_vld,
    l_TBlock_1_1_2_0153_out,
    l_TBlock_1_1_2_0153_out_ap_vld,
    l_TBlock_1_1_1_0152_out,
    l_TBlock_1_1_1_0152_out_ap_vld,
    l_TBlock_1_1_0_0151_out,
    l_TBlock_1_1_0_0151_out_ap_vld,
    l_TBlock_1_0_3_0150_out,
    l_TBlock_1_0_3_0150_out_ap_vld,
    l_TBlock_1_0_2_0149_out,
    l_TBlock_1_0_2_0149_out_ap_vld,
    l_TBlock_1_0_1_0148_out,
    l_TBlock_1_0_1_0148_out_ap_vld,
    l_TBlock_1_0_0_0147_out,
    l_TBlock_1_0_0_0147_out_ap_vld,
    l_TBlock_0_3_3_0146_out,
    l_TBlock_0_3_3_0146_out_ap_vld,
    l_TBlock_0_3_2_0145_out,
    l_TBlock_0_3_2_0145_out_ap_vld,
    l_TBlock_0_3_1_0144_out,
    l_TBlock_0_3_1_0144_out_ap_vld,
    l_TBlock_0_3_0_0143_out,
    l_TBlock_0_3_0_0143_out_ap_vld,
    l_TBlock_0_2_3_0142_out,
    l_TBlock_0_2_3_0142_out_ap_vld,
    l_TBlock_0_2_2_0141_out,
    l_TBlock_0_2_2_0141_out_ap_vld,
    l_TBlock_0_2_1_0140_out,
    l_TBlock_0_2_1_0140_out_ap_vld,
    l_TBlock_0_2_0_0139_out,
    l_TBlock_0_2_0_0139_out_ap_vld,
    l_TBlock_0_1_3_0138_out,
    l_TBlock_0_1_3_0138_out_ap_vld,
    l_TBlock_0_1_2_0137_out,
    l_TBlock_0_1_2_0137_out_ap_vld,
    l_TBlock_0_1_1_0136_out,
    l_TBlock_0_1_1_0136_out_ap_vld,
    l_TBlock_0_1_0_0135_out,
    l_TBlock_0_1_0_0135_out_ap_vld,
    l_TBlock_0_0_3_0134_out,
    l_TBlock_0_0_3_0134_out_ap_vld,
    l_TBlock_0_0_2_0133_out,
    l_TBlock_0_0_2_0133_out_ap_vld,
    l_TBlock_0_0_1_0132_out,
    l_TBlock_0_0_1_0132_out_ap_vld,
    l_TBlock_0_0_0_0131_out,
    l_TBlock_0_0_0_0131_out_ap_vld,
    l_TColl_0_0_0_constprop,
    l_TColl_0_0_0_constprop_ap_vld,
    l_TColl_0_1_0_constprop,
    l_TColl_0_1_0_constprop_ap_vld,
    l_TColl_0_2_0_constprop,
    l_TColl_0_2_0_constprop_ap_vld,
    l_TColl_0_3_0_constprop,
    l_TColl_0_3_0_constprop_ap_vld,
    l_TColl_1_0_0_constprop,
    l_TColl_1_0_0_constprop_ap_vld,
    l_TColl_1_1_0_constprop,
    l_TColl_1_1_0_constprop_ap_vld,
    l_TColl_1_2_0_constprop,
    l_TColl_1_2_0_constprop_ap_vld,
    l_TColl_1_3_0_constprop,
    l_TColl_1_3_0_constprop_ap_vld,
    l_TColl_2_0_0_constprop,
    l_TColl_2_0_0_constprop_ap_vld,
    l_TColl_2_1_0_constprop,
    l_TColl_2_1_0_constprop_ap_vld,
    l_TColl_2_2_0_constprop,
    l_TColl_2_2_0_constprop_ap_vld,
    l_TColl_2_3_0_constprop,
    l_TColl_2_3_0_constprop_ap_vld,
    l_TColl_0_0_1_constprop,
    l_TColl_0_0_1_constprop_ap_vld,
    l_TColl_0_1_1_constprop,
    l_TColl_0_1_1_constprop_ap_vld,
    l_TColl_0_2_1_constprop,
    l_TColl_0_2_1_constprop_ap_vld,
    l_TColl_0_3_1_constprop,
    l_TColl_0_3_1_constprop_ap_vld,
    l_TColl_1_0_1_constprop,
    l_TColl_1_0_1_constprop_ap_vld,
    l_TColl_1_1_1_constprop,
    l_TColl_1_1_1_constprop_ap_vld,
    l_TColl_1_2_1_constprop,
    l_TColl_1_2_1_constprop_ap_vld,
    l_TColl_1_3_1_constprop,
    l_TColl_1_3_1_constprop_ap_vld,
    l_TColl_2_0_1_constprop,
    l_TColl_2_0_1_constprop_ap_vld,
    l_TColl_2_1_1_constprop,
    l_TColl_2_1_1_constprop_ap_vld,
    l_TColl_2_2_1_constprop,
    l_TColl_2_2_1_constprop_ap_vld,
    l_TColl_2_3_1_constprop,
    l_TColl_2_3_1_constprop_ap_vld,
    l_TColl_0_0_2_constprop,
    l_TColl_0_0_2_constprop_ap_vld,
    l_TColl_0_1_2_constprop,
    l_TColl_0_1_2_constprop_ap_vld,
    l_TColl_0_2_2_constprop,
    l_TColl_0_2_2_constprop_ap_vld,
    l_TColl_0_3_2_constprop,
    l_TColl_0_3_2_constprop_ap_vld,
    l_TColl_1_0_2_constprop,
    l_TColl_1_0_2_constprop_ap_vld,
    l_TColl_1_1_2_constprop,
    l_TColl_1_1_2_constprop_ap_vld,
    l_TColl_1_2_2_constprop,
    l_TColl_1_2_2_constprop_ap_vld,
    l_TColl_1_3_2_constprop,
    l_TColl_1_3_2_constprop_ap_vld,
    l_TColl_2_0_2_constprop,
    l_TColl_2_0_2_constprop_ap_vld,
    l_TColl_2_1_2_constprop,
    l_TColl_2_1_2_constprop_ap_vld,
    l_TColl_2_2_2_constprop,
    l_TColl_2_2_2_constprop_ap_vld,
    l_TColl_2_3_2_constprop,
    l_TColl_2_3_2_constprop_ap_vld,
    l_TColl_0_0_3_constprop,
    l_TColl_0_0_3_constprop_ap_vld,
    l_TColl_0_1_3_constprop,
    l_TColl_0_1_3_constprop_ap_vld,
    l_TColl_0_2_3_constprop,
    l_TColl_0_2_3_constprop_ap_vld,
    l_TColl_0_3_3_constprop,
    l_TColl_0_3_3_constprop_ap_vld,
    l_TColl_1_0_3_constprop,
    l_TColl_1_0_3_constprop_ap_vld,
    l_TColl_1_1_3_constprop,
    l_TColl_1_1_3_constprop_ap_vld,
    l_TColl_1_2_3_constprop,
    l_TColl_1_2_3_constprop_ap_vld,
    l_TColl_1_3_3_constprop,
    l_TColl_1_3_3_constprop_ap_vld,
    l_TColl_2_0_3_constprop,
    l_TColl_2_0_3_constprop_ap_vld,
    l_TColl_2_1_3_constprop,
    l_TColl_2_1_3_constprop_ap_vld,
    l_TColl_2_2_3_constprop,
    l_TColl_2_2_3_constprop_ap_vld,
    l_TColl_2_3_3_constprop,
    l_TColl_2_3_3_constprop_ap_vld
);

    parameter ap_ST_fsm_pp0_stage0 = 78'd1;
    parameter ap_ST_fsm_pp0_stage1 = 78'd2;
    parameter ap_ST_fsm_pp0_stage2 = 78'd4;
    parameter ap_ST_fsm_pp0_stage3 = 78'd8;
    parameter ap_ST_fsm_pp0_stage4 = 78'd16;
    parameter ap_ST_fsm_pp0_stage5 = 78'd32;
    parameter ap_ST_fsm_pp0_stage6 = 78'd64;
    parameter ap_ST_fsm_pp0_stage7 = 78'd128;
    parameter ap_ST_fsm_pp0_stage8 = 78'd256;
    parameter ap_ST_fsm_pp0_stage9 = 78'd512;
    parameter ap_ST_fsm_pp0_stage10 = 78'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 78'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 78'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 78'd8192;
    parameter ap_ST_fsm_pp0_stage14 = 78'd16384;
    parameter ap_ST_fsm_pp0_stage15 = 78'd32768;
    parameter ap_ST_fsm_pp0_stage16 = 78'd65536;
    parameter ap_ST_fsm_pp0_stage17 = 78'd131072;
    parameter ap_ST_fsm_pp0_stage18 = 78'd262144;
    parameter ap_ST_fsm_pp0_stage19 = 78'd524288;
    parameter ap_ST_fsm_pp0_stage20 = 78'd1048576;
    parameter ap_ST_fsm_pp0_stage21 = 78'd2097152;
    parameter ap_ST_fsm_pp0_stage22 = 78'd4194304;
    parameter ap_ST_fsm_pp0_stage23 = 78'd8388608;
    parameter ap_ST_fsm_pp0_stage24 = 78'd16777216;
    parameter ap_ST_fsm_pp0_stage25 = 78'd33554432;
    parameter ap_ST_fsm_pp0_stage26 = 78'd67108864;
    parameter ap_ST_fsm_pp0_stage27 = 78'd134217728;
    parameter ap_ST_fsm_pp0_stage28 = 78'd268435456;
    parameter ap_ST_fsm_pp0_stage29 = 78'd536870912;
    parameter ap_ST_fsm_pp0_stage30 = 78'd1073741824;
    parameter ap_ST_fsm_pp0_stage31 = 78'd2147483648;
    parameter ap_ST_fsm_pp0_stage32 = 78'd4294967296;
    parameter ap_ST_fsm_pp0_stage33 = 78'd8589934592;
    parameter ap_ST_fsm_pp0_stage34 = 78'd17179869184;
    parameter ap_ST_fsm_pp0_stage35 = 78'd34359738368;
    parameter ap_ST_fsm_pp0_stage36 = 78'd68719476736;
    parameter ap_ST_fsm_pp0_stage37 = 78'd137438953472;
    parameter ap_ST_fsm_pp0_stage38 = 78'd274877906944;
    parameter ap_ST_fsm_pp0_stage39 = 78'd549755813888;
    parameter ap_ST_fsm_pp0_stage40 = 78'd1099511627776;
    parameter ap_ST_fsm_pp0_stage41 = 78'd2199023255552;
    parameter ap_ST_fsm_pp0_stage42 = 78'd4398046511104;
    parameter ap_ST_fsm_pp0_stage43 = 78'd8796093022208;
    parameter ap_ST_fsm_pp0_stage44 = 78'd17592186044416;
    parameter ap_ST_fsm_pp0_stage45 = 78'd35184372088832;
    parameter ap_ST_fsm_pp0_stage46 = 78'd70368744177664;
    parameter ap_ST_fsm_pp0_stage47 = 78'd140737488355328;
    parameter ap_ST_fsm_pp0_stage48 = 78'd281474976710656;
    parameter ap_ST_fsm_pp0_stage49 = 78'd562949953421312;
    parameter ap_ST_fsm_pp0_stage50 = 78'd1125899906842624;
    parameter ap_ST_fsm_pp0_stage51 = 78'd2251799813685248;
    parameter ap_ST_fsm_pp0_stage52 = 78'd4503599627370496;
    parameter ap_ST_fsm_pp0_stage53 = 78'd9007199254740992;
    parameter ap_ST_fsm_pp0_stage54 = 78'd18014398509481984;
    parameter ap_ST_fsm_pp0_stage55 = 78'd36028797018963968;
    parameter ap_ST_fsm_pp0_stage56 = 78'd72057594037927936;
    parameter ap_ST_fsm_pp0_stage57 = 78'd144115188075855872;
    parameter ap_ST_fsm_pp0_stage58 = 78'd288230376151711744;
    parameter ap_ST_fsm_pp0_stage59 = 78'd576460752303423488;
    parameter ap_ST_fsm_pp0_stage60 = 78'd1152921504606846976;
    parameter ap_ST_fsm_pp0_stage61 = 78'd2305843009213693952;
    parameter ap_ST_fsm_pp0_stage62 = 78'd4611686018427387904;
    parameter ap_ST_fsm_pp0_stage63 = 78'd9223372036854775808;
    parameter ap_ST_fsm_pp0_stage64 = 78'd18446744073709551616;
    parameter ap_ST_fsm_pp0_stage65 = 78'd36893488147419103232;
    parameter ap_ST_fsm_pp0_stage66 = 78'd73786976294838206464;
    parameter ap_ST_fsm_pp0_stage67 = 78'd147573952589676412928;
    parameter ap_ST_fsm_pp0_stage68 = 78'd295147905179352825856;
    parameter ap_ST_fsm_pp0_stage69 = 78'd590295810358705651712;
    parameter ap_ST_fsm_pp0_stage70 = 78'd1180591620717411303424;
    parameter ap_ST_fsm_pp0_stage71 = 78'd2361183241434822606848;
    parameter ap_ST_fsm_pp0_stage72 = 78'd4722366482869645213696;
    parameter ap_ST_fsm_pp0_stage73 = 78'd9444732965739290427392;
    parameter ap_ST_fsm_pp0_stage74 = 78'd18889465931478580854784;
    parameter ap_ST_fsm_pp0_stage75 = 78'd37778931862957161709568;
    parameter ap_ST_fsm_pp0_stage76 = 78'd75557863725914323419136;
    parameter ap_ST_fsm_pp0_stage77 = 78'd151115727451828646838272;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [63:0] l_TBlock_3_3_3_0194_out;
    output l_TBlock_3_3_3_0194_out_ap_vld;
    output [63:0] l_TBlock_3_3_2_0193_out;
    output l_TBlock_3_3_2_0193_out_ap_vld;
    output [63:0] l_TBlock_3_3_1_0192_out;
    output l_TBlock_3_3_1_0192_out_ap_vld;
    output [63:0] l_TBlock_3_3_0_0191_out;
    output l_TBlock_3_3_0_0191_out_ap_vld;
    output [63:0] l_TBlock_3_2_3_0190_out;
    output l_TBlock_3_2_3_0190_out_ap_vld;
    output [63:0] l_TBlock_3_2_2_0189_out;
    output l_TBlock_3_2_2_0189_out_ap_vld;
    output [63:0] l_TBlock_3_2_1_0188_out;
    output l_TBlock_3_2_1_0188_out_ap_vld;
    output [63:0] l_TBlock_3_2_0_0187_out;
    output l_TBlock_3_2_0_0187_out_ap_vld;
    output [63:0] l_TBlock_3_1_3_0186_out;
    output l_TBlock_3_1_3_0186_out_ap_vld;
    output [63:0] l_TBlock_3_1_2_0185_out;
    output l_TBlock_3_1_2_0185_out_ap_vld;
    output [63:0] l_TBlock_3_1_1_0184_out;
    output l_TBlock_3_1_1_0184_out_ap_vld;
    output [63:0] l_TBlock_3_1_0_0183_out;
    output l_TBlock_3_1_0_0183_out_ap_vld;
    output [63:0] l_TBlock_3_0_3_0182_out;
    output l_TBlock_3_0_3_0182_out_ap_vld;
    output [63:0] l_TBlock_3_0_2_0181_out;
    output l_TBlock_3_0_2_0181_out_ap_vld;
    output [63:0] l_TBlock_3_0_1_0180_out;
    output l_TBlock_3_0_1_0180_out_ap_vld;
    output [63:0] l_TBlock_3_0_0_0179_out;
    output l_TBlock_3_0_0_0179_out_ap_vld;
    output [63:0] l_TBlock_2_3_3_0178_out;
    output l_TBlock_2_3_3_0178_out_ap_vld;
    output [63:0] l_TBlock_2_3_2_0177_out;
    output l_TBlock_2_3_2_0177_out_ap_vld;
    output [63:0] l_TBlock_2_3_1_0176_out;
    output l_TBlock_2_3_1_0176_out_ap_vld;
    output [63:0] l_TBlock_2_3_0_0175_out;
    output l_TBlock_2_3_0_0175_out_ap_vld;
    output [63:0] l_TBlock_2_2_3_0174_out;
    output l_TBlock_2_2_3_0174_out_ap_vld;
    output [63:0] l_TBlock_2_2_2_0173_out;
    output l_TBlock_2_2_2_0173_out_ap_vld;
    output [63:0] l_TBlock_2_2_1_0172_out;
    output l_TBlock_2_2_1_0172_out_ap_vld;
    output [63:0] l_TBlock_2_2_0_0171_out;
    output l_TBlock_2_2_0_0171_out_ap_vld;
    output [63:0] l_TBlock_2_1_3_0170_out;
    output l_TBlock_2_1_3_0170_out_ap_vld;
    output [63:0] l_TBlock_2_1_2_0169_out;
    output l_TBlock_2_1_2_0169_out_ap_vld;
    output [63:0] l_TBlock_2_1_1_0168_out;
    output l_TBlock_2_1_1_0168_out_ap_vld;
    output [63:0] l_TBlock_2_1_0_0167_out;
    output l_TBlock_2_1_0_0167_out_ap_vld;
    output [63:0] l_TBlock_2_0_3_0166_out;
    output l_TBlock_2_0_3_0166_out_ap_vld;
    output [63:0] l_TBlock_2_0_2_0165_out;
    output l_TBlock_2_0_2_0165_out_ap_vld;
    output [63:0] l_TBlock_2_0_1_0164_out;
    output l_TBlock_2_0_1_0164_out_ap_vld;
    output [63:0] l_TBlock_2_0_0_0163_out;
    output l_TBlock_2_0_0_0163_out_ap_vld;
    output [63:0] l_TBlock_1_3_3_0162_out;
    output l_TBlock_1_3_3_0162_out_ap_vld;
    output [63:0] l_TBlock_1_3_2_0161_out;
    output l_TBlock_1_3_2_0161_out_ap_vld;
    output [63:0] l_TBlock_1_3_1_0160_out;
    output l_TBlock_1_3_1_0160_out_ap_vld;
    output [63:0] l_TBlock_1_3_0_0159_out;
    output l_TBlock_1_3_0_0159_out_ap_vld;
    output [63:0] l_TBlock_1_2_3_0158_out;
    output l_TBlock_1_2_3_0158_out_ap_vld;
    output [63:0] l_TBlock_1_2_2_0157_out;
    output l_TBlock_1_2_2_0157_out_ap_vld;
    output [63:0] l_TBlock_1_2_1_0156_out;
    output l_TBlock_1_2_1_0156_out_ap_vld;
    output [63:0] l_TBlock_1_2_0_0155_out;
    output l_TBlock_1_2_0_0155_out_ap_vld;
    output [63:0] l_TBlock_1_1_3_0154_out;
    output l_TBlock_1_1_3_0154_out_ap_vld;
    output [63:0] l_TBlock_1_1_2_0153_out;
    output l_TBlock_1_1_2_0153_out_ap_vld;
    output [63:0] l_TBlock_1_1_1_0152_out;
    output l_TBlock_1_1_1_0152_out_ap_vld;
    output [63:0] l_TBlock_1_1_0_0151_out;
    output l_TBlock_1_1_0_0151_out_ap_vld;
    output [63:0] l_TBlock_1_0_3_0150_out;
    output l_TBlock_1_0_3_0150_out_ap_vld;
    output [63:0] l_TBlock_1_0_2_0149_out;
    output l_TBlock_1_0_2_0149_out_ap_vld;
    output [63:0] l_TBlock_1_0_1_0148_out;
    output l_TBlock_1_0_1_0148_out_ap_vld;
    output [63:0] l_TBlock_1_0_0_0147_out;
    output l_TBlock_1_0_0_0147_out_ap_vld;
    output [63:0] l_TBlock_0_3_3_0146_out;
    output l_TBlock_0_3_3_0146_out_ap_vld;
    output [63:0] l_TBlock_0_3_2_0145_out;
    output l_TBlock_0_3_2_0145_out_ap_vld;
    output [63:0] l_TBlock_0_3_1_0144_out;
    output l_TBlock_0_3_1_0144_out_ap_vld;
    output [63:0] l_TBlock_0_3_0_0143_out;
    output l_TBlock_0_3_0_0143_out_ap_vld;
    output [63:0] l_TBlock_0_2_3_0142_out;
    output l_TBlock_0_2_3_0142_out_ap_vld;
    output [63:0] l_TBlock_0_2_2_0141_out;
    output l_TBlock_0_2_2_0141_out_ap_vld;
    output [63:0] l_TBlock_0_2_1_0140_out;
    output l_TBlock_0_2_1_0140_out_ap_vld;
    output [63:0] l_TBlock_0_2_0_0139_out;
    output l_TBlock_0_2_0_0139_out_ap_vld;
    output [63:0] l_TBlock_0_1_3_0138_out;
    output l_TBlock_0_1_3_0138_out_ap_vld;
    output [63:0] l_TBlock_0_1_2_0137_out;
    output l_TBlock_0_1_2_0137_out_ap_vld;
    output [63:0] l_TBlock_0_1_1_0136_out;
    output l_TBlock_0_1_1_0136_out_ap_vld;
    output [63:0] l_TBlock_0_1_0_0135_out;
    output l_TBlock_0_1_0_0135_out_ap_vld;
    output [63:0] l_TBlock_0_0_3_0134_out;
    output l_TBlock_0_0_3_0134_out_ap_vld;
    output [63:0] l_TBlock_0_0_2_0133_out;
    output l_TBlock_0_0_2_0133_out_ap_vld;
    output [63:0] l_TBlock_0_0_1_0132_out;
    output l_TBlock_0_0_1_0132_out_ap_vld;
    output [63:0] l_TBlock_0_0_0_0131_out;
    output l_TBlock_0_0_0_0131_out_ap_vld;
    output [63:0] l_TColl_0_0_0_constprop;
    output l_TColl_0_0_0_constprop_ap_vld;
    output [63:0] l_TColl_0_1_0_constprop;
    output l_TColl_0_1_0_constprop_ap_vld;
    output [63:0] l_TColl_0_2_0_constprop;
    output l_TColl_0_2_0_constprop_ap_vld;
    output [63:0] l_TColl_0_3_0_constprop;
    output l_TColl_0_3_0_constprop_ap_vld;
    output [63:0] l_TColl_1_0_0_constprop;
    output l_TColl_1_0_0_constprop_ap_vld;
    output [63:0] l_TColl_1_1_0_constprop;
    output l_TColl_1_1_0_constprop_ap_vld;
    output [63:0] l_TColl_1_2_0_constprop;
    output l_TColl_1_2_0_constprop_ap_vld;
    output [63:0] l_TColl_1_3_0_constprop;
    output l_TColl_1_3_0_constprop_ap_vld;
    output [63:0] l_TColl_2_0_0_constprop;
    output l_TColl_2_0_0_constprop_ap_vld;
    output [63:0] l_TColl_2_1_0_constprop;
    output l_TColl_2_1_0_constprop_ap_vld;
    output [63:0] l_TColl_2_2_0_constprop;
    output l_TColl_2_2_0_constprop_ap_vld;
    output [63:0] l_TColl_2_3_0_constprop;
    output l_TColl_2_3_0_constprop_ap_vld;
    output [63:0] l_TColl_0_0_1_constprop;
    output l_TColl_0_0_1_constprop_ap_vld;
    output [63:0] l_TColl_0_1_1_constprop;
    output l_TColl_0_1_1_constprop_ap_vld;
    output [63:0] l_TColl_0_2_1_constprop;
    output l_TColl_0_2_1_constprop_ap_vld;
    output [63:0] l_TColl_0_3_1_constprop;
    output l_TColl_0_3_1_constprop_ap_vld;
    output [63:0] l_TColl_1_0_1_constprop;
    output l_TColl_1_0_1_constprop_ap_vld;
    output [63:0] l_TColl_1_1_1_constprop;
    output l_TColl_1_1_1_constprop_ap_vld;
    output [63:0] l_TColl_1_2_1_constprop;
    output l_TColl_1_2_1_constprop_ap_vld;
    output [63:0] l_TColl_1_3_1_constprop;
    output l_TColl_1_3_1_constprop_ap_vld;
    output [63:0] l_TColl_2_0_1_constprop;
    output l_TColl_2_0_1_constprop_ap_vld;
    output [63:0] l_TColl_2_1_1_constprop;
    output l_TColl_2_1_1_constprop_ap_vld;
    output [63:0] l_TColl_2_2_1_constprop;
    output l_TColl_2_2_1_constprop_ap_vld;
    output [63:0] l_TColl_2_3_1_constprop;
    output l_TColl_2_3_1_constprop_ap_vld;
    output [63:0] l_TColl_0_0_2_constprop;
    output l_TColl_0_0_2_constprop_ap_vld;
    output [63:0] l_TColl_0_1_2_constprop;
    output l_TColl_0_1_2_constprop_ap_vld;
    output [63:0] l_TColl_0_2_2_constprop;
    output l_TColl_0_2_2_constprop_ap_vld;
    output [63:0] l_TColl_0_3_2_constprop;
    output l_TColl_0_3_2_constprop_ap_vld;
    output [63:0] l_TColl_1_0_2_constprop;
    output l_TColl_1_0_2_constprop_ap_vld;
    output [63:0] l_TColl_1_1_2_constprop;
    output l_TColl_1_1_2_constprop_ap_vld;
    output [63:0] l_TColl_1_2_2_constprop;
    output l_TColl_1_2_2_constprop_ap_vld;
    output [63:0] l_TColl_1_3_2_constprop;
    output l_TColl_1_3_2_constprop_ap_vld;
    output [63:0] l_TColl_2_0_2_constprop;
    output l_TColl_2_0_2_constprop_ap_vld;
    output [63:0] l_TColl_2_1_2_constprop;
    output l_TColl_2_1_2_constprop_ap_vld;
    output [63:0] l_TColl_2_2_2_constprop;
    output l_TColl_2_2_2_constprop_ap_vld;
    output [63:0] l_TColl_2_3_2_constprop;
    output l_TColl_2_3_2_constprop_ap_vld;
    output [63:0] l_TColl_0_0_3_constprop;
    output l_TColl_0_0_3_constprop_ap_vld;
    output [63:0] l_TColl_0_1_3_constprop;
    output l_TColl_0_1_3_constprop_ap_vld;
    output [63:0] l_TColl_0_2_3_constprop;
    output l_TColl_0_2_3_constprop_ap_vld;
    output [63:0] l_TColl_0_3_3_constprop;
    output l_TColl_0_3_3_constprop_ap_vld;
    output [63:0] l_TColl_1_0_3_constprop;
    output l_TColl_1_0_3_constprop_ap_vld;
    output [63:0] l_TColl_1_1_3_constprop;
    output l_TColl_1_1_3_constprop_ap_vld;
    output [63:0] l_TColl_1_2_3_constprop;
    output l_TColl_1_2_3_constprop_ap_vld;
    output [63:0] l_TColl_1_3_3_constprop;
    output l_TColl_1_3_3_constprop_ap_vld;
    output [63:0] l_TColl_2_0_3_constprop;
    output l_TColl_2_0_3_constprop_ap_vld;
    output [63:0] l_TColl_2_1_3_constprop;
    output l_TColl_2_1_3_constprop_ap_vld;
    output [63:0] l_TColl_2_2_3_constprop;
    output l_TColl_2_2_3_constprop_ap_vld;
    output [63:0] l_TColl_2_3_3_constprop;
    output l_TColl_2_3_3_constprop_ap_vld;

    reg ap_idle;
    reg l_TBlock_3_3_3_0194_out_ap_vld;
    reg l_TBlock_3_3_2_0193_out_ap_vld;
    reg l_TBlock_3_3_1_0192_out_ap_vld;
    reg l_TBlock_3_3_0_0191_out_ap_vld;
    reg l_TBlock_3_2_3_0190_out_ap_vld;
    reg l_TBlock_3_2_2_0189_out_ap_vld;
    reg l_TBlock_3_2_1_0188_out_ap_vld;
    reg l_TBlock_3_2_0_0187_out_ap_vld;
    reg l_TBlock_3_1_3_0186_out_ap_vld;
    reg l_TBlock_3_1_2_0185_out_ap_vld;
    reg l_TBlock_3_1_1_0184_out_ap_vld;
    reg l_TBlock_3_1_0_0183_out_ap_vld;
    reg l_TBlock_3_0_3_0182_out_ap_vld;
    reg l_TBlock_3_0_2_0181_out_ap_vld;
    reg l_TBlock_3_0_1_0180_out_ap_vld;
    reg l_TBlock_3_0_0_0179_out_ap_vld;
    reg l_TBlock_2_3_3_0178_out_ap_vld;
    reg l_TBlock_2_3_2_0177_out_ap_vld;
    reg l_TBlock_2_3_1_0176_out_ap_vld;
    reg l_TBlock_2_3_0_0175_out_ap_vld;
    reg l_TBlock_2_2_3_0174_out_ap_vld;
    reg l_TBlock_2_2_2_0173_out_ap_vld;
    reg l_TBlock_2_2_1_0172_out_ap_vld;
    reg l_TBlock_2_2_0_0171_out_ap_vld;
    reg l_TBlock_2_1_3_0170_out_ap_vld;
    reg l_TBlock_2_1_2_0169_out_ap_vld;
    reg l_TBlock_2_1_1_0168_out_ap_vld;
    reg l_TBlock_2_1_0_0167_out_ap_vld;
    reg l_TBlock_2_0_3_0166_out_ap_vld;
    reg l_TBlock_2_0_2_0165_out_ap_vld;
    reg l_TBlock_2_0_1_0164_out_ap_vld;
    reg l_TBlock_2_0_0_0163_out_ap_vld;
    reg l_TBlock_1_3_3_0162_out_ap_vld;
    reg l_TBlock_1_3_2_0161_out_ap_vld;
    reg l_TBlock_1_3_1_0160_out_ap_vld;
    reg l_TBlock_1_3_0_0159_out_ap_vld;
    reg l_TBlock_1_2_3_0158_out_ap_vld;
    reg l_TBlock_1_2_2_0157_out_ap_vld;
    reg l_TBlock_1_2_1_0156_out_ap_vld;
    reg l_TBlock_1_2_0_0155_out_ap_vld;
    reg l_TBlock_1_1_3_0154_out_ap_vld;
    reg l_TBlock_1_1_2_0153_out_ap_vld;
    reg l_TBlock_1_1_1_0152_out_ap_vld;
    reg l_TBlock_1_1_0_0151_out_ap_vld;
    reg l_TBlock_1_0_3_0150_out_ap_vld;
    reg l_TBlock_1_0_2_0149_out_ap_vld;
    reg l_TBlock_1_0_1_0148_out_ap_vld;
    reg l_TBlock_1_0_0_0147_out_ap_vld;
    reg l_TBlock_0_3_3_0146_out_ap_vld;
    reg l_TBlock_0_3_2_0145_out_ap_vld;
    reg l_TBlock_0_3_1_0144_out_ap_vld;
    reg l_TBlock_0_3_0_0143_out_ap_vld;
    reg l_TBlock_0_2_3_0142_out_ap_vld;
    reg l_TBlock_0_2_2_0141_out_ap_vld;
    reg l_TBlock_0_2_1_0140_out_ap_vld;
    reg l_TBlock_0_2_0_0139_out_ap_vld;
    reg l_TBlock_0_1_3_0138_out_ap_vld;
    reg l_TBlock_0_1_2_0137_out_ap_vld;
    reg l_TBlock_0_1_1_0136_out_ap_vld;
    reg l_TBlock_0_1_0_0135_out_ap_vld;
    reg l_TBlock_0_0_3_0134_out_ap_vld;
    reg l_TBlock_0_0_2_0133_out_ap_vld;
    reg l_TBlock_0_0_1_0132_out_ap_vld;
    reg l_TBlock_0_0_0_0131_out_ap_vld;
    reg l_TColl_0_0_0_constprop_ap_vld;
    reg l_TColl_0_1_0_constprop_ap_vld;
    reg l_TColl_0_2_0_constprop_ap_vld;
    reg l_TColl_0_3_0_constprop_ap_vld;
    reg l_TColl_1_0_0_constprop_ap_vld;
    reg l_TColl_1_1_0_constprop_ap_vld;
    reg l_TColl_1_2_0_constprop_ap_vld;
    reg l_TColl_1_3_0_constprop_ap_vld;
    reg l_TColl_2_0_0_constprop_ap_vld;
    reg l_TColl_2_1_0_constprop_ap_vld;
    reg l_TColl_2_2_0_constprop_ap_vld;
    reg l_TColl_2_3_0_constprop_ap_vld;
    reg l_TColl_0_0_1_constprop_ap_vld;
    reg l_TColl_0_1_1_constprop_ap_vld;
    reg l_TColl_0_2_1_constprop_ap_vld;
    reg l_TColl_0_3_1_constprop_ap_vld;
    reg l_TColl_1_0_1_constprop_ap_vld;
    reg l_TColl_1_1_1_constprop_ap_vld;
    reg l_TColl_1_2_1_constprop_ap_vld;
    reg l_TColl_1_3_1_constprop_ap_vld;
    reg l_TColl_2_0_1_constprop_ap_vld;
    reg l_TColl_2_1_1_constprop_ap_vld;
    reg l_TColl_2_2_1_constprop_ap_vld;
    reg l_TColl_2_3_1_constprop_ap_vld;
    reg l_TColl_0_0_2_constprop_ap_vld;
    reg l_TColl_0_1_2_constprop_ap_vld;
    reg l_TColl_0_2_2_constprop_ap_vld;
    reg l_TColl_0_3_2_constprop_ap_vld;
    reg l_TColl_1_0_2_constprop_ap_vld;
    reg l_TColl_1_1_2_constprop_ap_vld;
    reg l_TColl_1_2_2_constprop_ap_vld;
    reg l_TColl_1_3_2_constprop_ap_vld;
    reg l_TColl_2_0_2_constprop_ap_vld;
    reg l_TColl_2_1_2_constprop_ap_vld;
    reg l_TColl_2_2_2_constprop_ap_vld;
    reg l_TColl_2_3_2_constprop_ap_vld;
    reg l_TColl_0_0_3_constprop_ap_vld;
    reg l_TColl_0_1_3_constprop_ap_vld;
    reg l_TColl_0_2_3_constprop_ap_vld;
    reg l_TColl_0_3_3_constprop_ap_vld;
    reg l_TColl_1_0_3_constprop_ap_vld;
    reg l_TColl_1_1_3_constprop_ap_vld;
    reg l_TColl_1_2_3_constprop_ap_vld;
    reg l_TColl_1_3_3_constprop_ap_vld;
    reg l_TColl_2_0_3_constprop_ap_vld;
    reg l_TColl_2_1_3_constprop_ap_vld;
    reg l_TColl_2_2_3_constprop_ap_vld;
    reg l_TColl_2_3_3_constprop_ap_vld;

    (* fsm_encoding = "none" *) reg   [77:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_subdone;
    reg   [0:0] icmp_ln69_reg_2958;
    reg    ap_condition_exit_pp0_iter0_stage1;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_CS_fsm_pp0_stage77;
    wire    ap_block_pp0_stage77_subdone;
    wire    ap_block_pp0_stage0_11001;
    wire   [0:0] icmp_ln69_fu_1064_p2;
    wire   [1:0] trunc_ln69_fu_1076_p1;
    reg   [1:0] trunc_ln69_reg_2962;
    wire   [63:0] tmp_fu_1080_p6;
    reg   [63:0] tmp_reg_2967;
    wire   [63:0] tmp_s_fu_1094_p6;
    reg   [63:0] tmp_s_reg_2972;
    wire   [63:0] tmp_270_fu_1108_p6;
    reg   [63:0] tmp_270_reg_2977;
    wire    ap_block_pp0_stage1_11001;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_0;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_1;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_2;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_3;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_4;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_5;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_6;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_7;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_8;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_9;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_10;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_11;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_12;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_13;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_14;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_15;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_16;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_17;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_18;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_19;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_20;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_21;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_22;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_23;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_24;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_25;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_26;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_27;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_28;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_29;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_30;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_31;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_32;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_33;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_34;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_35;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_36;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_37;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_38;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_39;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_40;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_41;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_42;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_43;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_44;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_45;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_46;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_47;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_48;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_49;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_50;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_51;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_52;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_53;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_54;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_55;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_56;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_57;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_58;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_59;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_60;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_61;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_62;
    wire   [63:0] grp_rpyxyzToH_double_s_fu_984_ap_return_63;
    wire    ap_block_pp0_stage1;
    wire    ap_block_pp0_stage0;
    reg   [2:0] i_1_fu_276;
    wire   [2:0] add_ln69_fu_1070_p2;
    wire    ap_loop_init;
    reg   [2:0] ap_sig_allocacmp_i;
    reg   [63:0] l_TBlock_0_0_0_0131_fu_280;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_0_0_0131_load_1;
    reg   [63:0] l_TBlock_0_0_1_0132_fu_284;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_0_1_0132_load_1;
    reg   [63:0] l_TBlock_0_0_2_0133_fu_288;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_0_2_0133_load_1;
    reg   [63:0] l_TBlock_0_0_3_0134_fu_292;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_0_3_0134_load_1;
    reg   [63:0] l_TBlock_0_1_0_0135_fu_296;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_1_0_0135_load_1;
    reg   [63:0] l_TBlock_0_1_1_0136_fu_300;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_1_1_0136_load_1;
    reg   [63:0] l_TBlock_0_1_2_0137_fu_304;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_1_2_0137_load_1;
    reg   [63:0] l_TBlock_0_1_3_0138_fu_308;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_1_3_0138_load_1;
    reg   [63:0] l_TBlock_0_2_0_0139_fu_312;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_2_0_0139_load_1;
    reg   [63:0] l_TBlock_0_2_1_0140_fu_316;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_2_1_0140_load_1;
    reg   [63:0] l_TBlock_0_2_2_0141_fu_320;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_2_2_0141_load_1;
    reg   [63:0] l_TBlock_0_2_3_0142_fu_324;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_2_3_0142_load_1;
    reg   [63:0] l_TBlock_0_3_0_0143_fu_328;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_3_0_0143_load_1;
    reg   [63:0] l_TBlock_0_3_1_0144_fu_332;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_3_1_0144_load_1;
    reg   [63:0] l_TBlock_0_3_2_0145_fu_336;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_3_2_0145_load_1;
    reg   [63:0] l_TBlock_0_3_3_0146_fu_340;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_0_3_3_0146_load_1;
    reg   [63:0] l_TBlock_1_0_0_0147_fu_344;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_0_0_0147_load_1;
    reg   [63:0] l_TBlock_1_0_1_0148_fu_348;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_0_1_0148_load_1;
    reg   [63:0] l_TBlock_1_0_2_0149_fu_352;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_0_2_0149_load_1;
    reg   [63:0] l_TBlock_1_0_3_0150_fu_356;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_0_3_0150_load_1;
    reg   [63:0] l_TBlock_1_1_0_0151_fu_360;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_1_0_0151_load_1;
    reg   [63:0] l_TBlock_1_1_1_0152_fu_364;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_1_1_0152_load_1;
    reg   [63:0] l_TBlock_1_1_2_0153_fu_368;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_1_2_0153_load_1;
    reg   [63:0] l_TBlock_1_1_3_0154_fu_372;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_1_3_0154_load_1;
    reg   [63:0] l_TBlock_1_2_0_0155_fu_376;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_2_0_0155_load_1;
    reg   [63:0] l_TBlock_1_2_1_0156_fu_380;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_2_1_0156_load_1;
    reg   [63:0] l_TBlock_1_2_2_0157_fu_384;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_2_2_0157_load_1;
    reg   [63:0] l_TBlock_1_2_3_0158_fu_388;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_2_3_0158_load_1;
    reg   [63:0] l_TBlock_1_3_0_0159_fu_392;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_3_0_0159_load_1;
    reg   [63:0] l_TBlock_1_3_1_0160_fu_396;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_3_1_0160_load_1;
    reg   [63:0] l_TBlock_1_3_2_0161_fu_400;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_3_2_0161_load_1;
    reg   [63:0] l_TBlock_1_3_3_0162_fu_404;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_1_3_3_0162_load_1;
    reg   [63:0] l_TBlock_2_0_0_0163_fu_408;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_0_0_0163_load_1;
    reg   [63:0] l_TBlock_2_0_1_0164_fu_412;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_0_1_0164_load_1;
    reg   [63:0] l_TBlock_2_0_2_0165_fu_416;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_0_2_0165_load_1;
    reg   [63:0] l_TBlock_2_0_3_0166_fu_420;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_0_3_0166_load_1;
    reg   [63:0] l_TBlock_2_1_0_0167_fu_424;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_1_0_0167_load_1;
    reg   [63:0] l_TBlock_2_1_1_0168_fu_428;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_1_1_0168_load_1;
    reg   [63:0] l_TBlock_2_1_2_0169_fu_432;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_1_2_0169_load_1;
    reg   [63:0] l_TBlock_2_1_3_0170_fu_436;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_1_3_0170_load_1;
    reg   [63:0] l_TBlock_2_2_0_0171_fu_440;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_2_0_0171_load_1;
    reg   [63:0] l_TBlock_2_2_1_0172_fu_444;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_2_1_0172_load_1;
    reg   [63:0] l_TBlock_2_2_2_0173_fu_448;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_2_2_0173_load_1;
    reg   [63:0] l_TBlock_2_2_3_0174_fu_452;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_2_3_0174_load_1;
    reg   [63:0] l_TBlock_2_3_0_0175_fu_456;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_3_0_0175_load_1;
    reg   [63:0] l_TBlock_2_3_1_0176_fu_460;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_3_1_0176_load_1;
    reg   [63:0] l_TBlock_2_3_2_0177_fu_464;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_3_2_0177_load_1;
    reg   [63:0] l_TBlock_2_3_3_0178_fu_468;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_2_3_3_0178_load_1;
    reg   [63:0] l_TBlock_3_0_0_0179_fu_472;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_0_0_0179_load_1;
    reg   [63:0] l_TBlock_3_0_1_0180_fu_476;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_0_1_0180_load_1;
    reg   [63:0] l_TBlock_3_0_2_0181_fu_480;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_0_2_0181_load_1;
    reg   [63:0] l_TBlock_3_0_3_0182_fu_484;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_0_3_0182_load_1;
    reg   [63:0] l_TBlock_3_1_0_0183_fu_488;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_1_0_0183_load_1;
    reg   [63:0] l_TBlock_3_1_1_0184_fu_492;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_1_1_0184_load_1;
    reg   [63:0] l_TBlock_3_1_2_0185_fu_496;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_1_2_0185_load_1;
    reg   [63:0] l_TBlock_3_1_3_0186_fu_500;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_1_3_0186_load_1;
    reg   [63:0] l_TBlock_3_2_0_0187_fu_504;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_2_0_0187_load_1;
    reg   [63:0] l_TBlock_3_2_1_0188_fu_508;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_2_1_0188_load_1;
    reg   [63:0] l_TBlock_3_2_2_0189_fu_512;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_2_2_0189_load_1;
    reg   [63:0] l_TBlock_3_2_3_0190_fu_516;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_2_3_0190_load_1;
    reg   [63:0] l_TBlock_3_3_0_0191_fu_520;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_3_0_0191_load_1;
    reg   [63:0] l_TBlock_3_3_1_0192_fu_524;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_3_1_0192_load_1;
    reg   [63:0] l_TBlock_3_3_2_0193_fu_528;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_3_2_0193_load_1;
    reg   [63:0] l_TBlock_3_3_3_0194_fu_532;
    reg   [63:0] ap_sig_allocacmp_l_TBlock_3_3_3_0194_load_1;
    wire    ap_block_pp0_stage1_01001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [77:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to1;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    wire    ap_block_pp0_stage9_subdone;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_block_pp0_stage13_subdone;
    wire    ap_block_pp0_stage14_subdone;
    wire    ap_block_pp0_stage15_subdone;
    wire    ap_block_pp0_stage16_subdone;
    wire    ap_block_pp0_stage17_subdone;
    wire    ap_block_pp0_stage18_subdone;
    wire    ap_block_pp0_stage19_subdone;
    wire    ap_block_pp0_stage20_subdone;
    wire    ap_block_pp0_stage21_subdone;
    wire    ap_block_pp0_stage22_subdone;
    wire    ap_block_pp0_stage23_subdone;
    wire    ap_block_pp0_stage24_subdone;
    wire    ap_block_pp0_stage25_subdone;
    wire    ap_block_pp0_stage26_subdone;
    wire    ap_block_pp0_stage27_subdone;
    wire    ap_block_pp0_stage28_subdone;
    wire    ap_block_pp0_stage29_subdone;
    wire    ap_block_pp0_stage30_subdone;
    wire    ap_block_pp0_stage31_subdone;
    wire    ap_block_pp0_stage32_subdone;
    wire    ap_block_pp0_stage33_subdone;
    wire    ap_block_pp0_stage34_subdone;
    wire    ap_block_pp0_stage35_subdone;
    wire    ap_block_pp0_stage36_subdone;
    wire    ap_block_pp0_stage37_subdone;
    wire    ap_block_pp0_stage38_subdone;
    wire    ap_block_pp0_stage39_subdone;
    wire    ap_block_pp0_stage40_subdone;
    wire    ap_block_pp0_stage41_subdone;
    wire    ap_block_pp0_stage42_subdone;
    wire    ap_block_pp0_stage43_subdone;
    wire    ap_block_pp0_stage44_subdone;
    wire    ap_block_pp0_stage45_subdone;
    wire    ap_block_pp0_stage46_subdone;
    wire    ap_block_pp0_stage47_subdone;
    wire    ap_block_pp0_stage48_subdone;
    wire    ap_block_pp0_stage49_subdone;
    wire    ap_block_pp0_stage50_subdone;
    wire    ap_block_pp0_stage51_subdone;
    wire    ap_block_pp0_stage52_subdone;
    wire    ap_block_pp0_stage53_subdone;
    wire    ap_block_pp0_stage54_subdone;
    wire    ap_block_pp0_stage55_subdone;
    wire    ap_block_pp0_stage56_subdone;
    wire    ap_block_pp0_stage57_subdone;
    wire    ap_block_pp0_stage58_subdone;
    wire    ap_block_pp0_stage59_subdone;
    wire    ap_block_pp0_stage60_subdone;
    wire    ap_block_pp0_stage61_subdone;
    wire    ap_block_pp0_stage62_subdone;
    wire    ap_block_pp0_stage63_subdone;
    wire    ap_block_pp0_stage64_subdone;
    wire    ap_block_pp0_stage65_subdone;
    wire    ap_block_pp0_stage66_subdone;
    wire    ap_block_pp0_stage67_subdone;
    wire    ap_block_pp0_stage68_subdone;
    wire    ap_block_pp0_stage69_subdone;
    wire    ap_block_pp0_stage70_subdone;
    wire    ap_block_pp0_stage71_subdone;
    wire    ap_block_pp0_stage72_subdone;
    wire    ap_block_pp0_stage73_subdone;
    wire    ap_block_pp0_stage74_subdone;
    wire    ap_block_pp0_stage75_subdone;
    wire    ap_block_pp0_stage76_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 78'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 i_1_fu_276 = 3'd0;
        #0 l_TBlock_0_0_0_0131_fu_280 = 64'd0;
        #0 l_TBlock_0_0_1_0132_fu_284 = 64'd0;
        #0 l_TBlock_0_0_2_0133_fu_288 = 64'd0;
        #0 l_TBlock_0_0_3_0134_fu_292 = 64'd0;
        #0 l_TBlock_0_1_0_0135_fu_296 = 64'd0;
        #0 l_TBlock_0_1_1_0136_fu_300 = 64'd0;
        #0 l_TBlock_0_1_2_0137_fu_304 = 64'd0;
        #0 l_TBlock_0_1_3_0138_fu_308 = 64'd0;
        #0 l_TBlock_0_2_0_0139_fu_312 = 64'd0;
        #0 l_TBlock_0_2_1_0140_fu_316 = 64'd0;
        #0 l_TBlock_0_2_2_0141_fu_320 = 64'd0;
        #0 l_TBlock_0_2_3_0142_fu_324 = 64'd0;
        #0 l_TBlock_0_3_0_0143_fu_328 = 64'd0;
        #0 l_TBlock_0_3_1_0144_fu_332 = 64'd0;
        #0 l_TBlock_0_3_2_0145_fu_336 = 64'd0;
        #0 l_TBlock_0_3_3_0146_fu_340 = 64'd0;
        #0 l_TBlock_1_0_0_0147_fu_344 = 64'd0;
        #0 l_TBlock_1_0_1_0148_fu_348 = 64'd0;
        #0 l_TBlock_1_0_2_0149_fu_352 = 64'd0;
        #0 l_TBlock_1_0_3_0150_fu_356 = 64'd0;
        #0 l_TBlock_1_1_0_0151_fu_360 = 64'd0;
        #0 l_TBlock_1_1_1_0152_fu_364 = 64'd0;
        #0 l_TBlock_1_1_2_0153_fu_368 = 64'd0;
        #0 l_TBlock_1_1_3_0154_fu_372 = 64'd0;
        #0 l_TBlock_1_2_0_0155_fu_376 = 64'd0;
        #0 l_TBlock_1_2_1_0156_fu_380 = 64'd0;
        #0 l_TBlock_1_2_2_0157_fu_384 = 64'd0;
        #0 l_TBlock_1_2_3_0158_fu_388 = 64'd0;
        #0 l_TBlock_1_3_0_0159_fu_392 = 64'd0;
        #0 l_TBlock_1_3_1_0160_fu_396 = 64'd0;
        #0 l_TBlock_1_3_2_0161_fu_400 = 64'd0;
        #0 l_TBlock_1_3_3_0162_fu_404 = 64'd0;
        #0 l_TBlock_2_0_0_0163_fu_408 = 64'd0;
        #0 l_TBlock_2_0_1_0164_fu_412 = 64'd0;
        #0 l_TBlock_2_0_2_0165_fu_416 = 64'd0;
        #0 l_TBlock_2_0_3_0166_fu_420 = 64'd0;
        #0 l_TBlock_2_1_0_0167_fu_424 = 64'd0;
        #0 l_TBlock_2_1_1_0168_fu_428 = 64'd0;
        #0 l_TBlock_2_1_2_0169_fu_432 = 64'd0;
        #0 l_TBlock_2_1_3_0170_fu_436 = 64'd0;
        #0 l_TBlock_2_2_0_0171_fu_440 = 64'd0;
        #0 l_TBlock_2_2_1_0172_fu_444 = 64'd0;
        #0 l_TBlock_2_2_2_0173_fu_448 = 64'd0;
        #0 l_TBlock_2_2_3_0174_fu_452 = 64'd0;
        #0 l_TBlock_2_3_0_0175_fu_456 = 64'd0;
        #0 l_TBlock_2_3_1_0176_fu_460 = 64'd0;
        #0 l_TBlock_2_3_2_0177_fu_464 = 64'd0;
        #0 l_TBlock_2_3_3_0178_fu_468 = 64'd0;
        #0 l_TBlock_3_0_0_0179_fu_472 = 64'd0;
        #0 l_TBlock_3_0_1_0180_fu_476 = 64'd0;
        #0 l_TBlock_3_0_2_0181_fu_480 = 64'd0;
        #0 l_TBlock_3_0_3_0182_fu_484 = 64'd0;
        #0 l_TBlock_3_1_0_0183_fu_488 = 64'd0;
        #0 l_TBlock_3_1_1_0184_fu_492 = 64'd0;
        #0 l_TBlock_3_1_2_0185_fu_496 = 64'd0;
        #0 l_TBlock_3_1_3_0186_fu_500 = 64'd0;
        #0 l_TBlock_3_2_0_0187_fu_504 = 64'd0;
        #0 l_TBlock_3_2_1_0188_fu_508 = 64'd0;
        #0 l_TBlock_3_2_2_0189_fu_512 = 64'd0;
        #0 l_TBlock_3_2_3_0190_fu_516 = 64'd0;
        #0 l_TBlock_3_3_0_0191_fu_520 = 64'd0;
        #0 l_TBlock_3_3_1_0192_fu_524 = 64'd0;
        #0 l_TBlock_3_3_2_0193_fu_528 = 64'd0;
        #0 l_TBlock_3_3_3_0194_fu_532 = 64'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_rpyxyzToH_double_s grp_rpyxyzToH_double_s_fu_984 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .x(tmp_reg_2967),
        .y(tmp_s_reg_2972),
        .z(tmp_270_reg_2977),
        .p_read(ap_sig_allocacmp_l_TBlock_0_0_0_0131_load_1),
        .p_read1(ap_sig_allocacmp_l_TBlock_0_0_1_0132_load_1),
        .p_read2(ap_sig_allocacmp_l_TBlock_0_0_2_0133_load_1),
        .p_read3(ap_sig_allocacmp_l_TBlock_0_0_3_0134_load_1),
        .p_read4(ap_sig_allocacmp_l_TBlock_0_1_0_0135_load_1),
        .p_read5(ap_sig_allocacmp_l_TBlock_0_1_1_0136_load_1),
        .p_read6(ap_sig_allocacmp_l_TBlock_0_1_2_0137_load_1),
        .p_read7(ap_sig_allocacmp_l_TBlock_0_1_3_0138_load_1),
        .p_read8(ap_sig_allocacmp_l_TBlock_0_2_0_0139_load_1),
        .p_read9(ap_sig_allocacmp_l_TBlock_0_2_1_0140_load_1),
        .p_read10(ap_sig_allocacmp_l_TBlock_0_2_2_0141_load_1),
        .p_read11(ap_sig_allocacmp_l_TBlock_0_2_3_0142_load_1),
        .p_read12(ap_sig_allocacmp_l_TBlock_0_3_0_0143_load_1),
        .p_read13(ap_sig_allocacmp_l_TBlock_0_3_1_0144_load_1),
        .p_read14(ap_sig_allocacmp_l_TBlock_0_3_2_0145_load_1),
        .p_read15(ap_sig_allocacmp_l_TBlock_0_3_3_0146_load_1),
        .p_read16(ap_sig_allocacmp_l_TBlock_1_0_0_0147_load_1),
        .p_read17(ap_sig_allocacmp_l_TBlock_1_0_1_0148_load_1),
        .p_read18(ap_sig_allocacmp_l_TBlock_1_0_2_0149_load_1),
        .p_read19(ap_sig_allocacmp_l_TBlock_1_0_3_0150_load_1),
        .p_read20(ap_sig_allocacmp_l_TBlock_1_1_0_0151_load_1),
        .p_read21(ap_sig_allocacmp_l_TBlock_1_1_1_0152_load_1),
        .p_read22(ap_sig_allocacmp_l_TBlock_1_1_2_0153_load_1),
        .p_read23(ap_sig_allocacmp_l_TBlock_1_1_3_0154_load_1),
        .p_read24(ap_sig_allocacmp_l_TBlock_1_2_0_0155_load_1),
        .p_read25(ap_sig_allocacmp_l_TBlock_1_2_1_0156_load_1),
        .p_read26(ap_sig_allocacmp_l_TBlock_1_2_2_0157_load_1),
        .p_read27(ap_sig_allocacmp_l_TBlock_1_2_3_0158_load_1),
        .p_read28(ap_sig_allocacmp_l_TBlock_1_3_0_0159_load_1),
        .p_read29(ap_sig_allocacmp_l_TBlock_1_3_1_0160_load_1),
        .p_read30(ap_sig_allocacmp_l_TBlock_1_3_2_0161_load_1),
        .p_read31(ap_sig_allocacmp_l_TBlock_1_3_3_0162_load_1),
        .p_read32(ap_sig_allocacmp_l_TBlock_2_0_0_0163_load_1),
        .p_read33(ap_sig_allocacmp_l_TBlock_2_0_1_0164_load_1),
        .p_read34(ap_sig_allocacmp_l_TBlock_2_0_2_0165_load_1),
        .p_read35(ap_sig_allocacmp_l_TBlock_2_0_3_0166_load_1),
        .p_read36(ap_sig_allocacmp_l_TBlock_2_1_0_0167_load_1),
        .p_read37(ap_sig_allocacmp_l_TBlock_2_1_1_0168_load_1),
        .p_read38(ap_sig_allocacmp_l_TBlock_2_1_2_0169_load_1),
        .p_read39(ap_sig_allocacmp_l_TBlock_2_1_3_0170_load_1),
        .p_read40(ap_sig_allocacmp_l_TBlock_2_2_0_0171_load_1),
        .p_read41(ap_sig_allocacmp_l_TBlock_2_2_1_0172_load_1),
        .p_read42(ap_sig_allocacmp_l_TBlock_2_2_2_0173_load_1),
        .p_read43(ap_sig_allocacmp_l_TBlock_2_2_3_0174_load_1),
        .p_read44(ap_sig_allocacmp_l_TBlock_2_3_0_0175_load_1),
        .p_read45(ap_sig_allocacmp_l_TBlock_2_3_1_0176_load_1),
        .p_read46(ap_sig_allocacmp_l_TBlock_2_3_2_0177_load_1),
        .p_read47(ap_sig_allocacmp_l_TBlock_2_3_3_0178_load_1),
        .p_read48(ap_sig_allocacmp_l_TBlock_3_0_0_0179_load_1),
        .p_read49(ap_sig_allocacmp_l_TBlock_3_0_1_0180_load_1),
        .p_read50(ap_sig_allocacmp_l_TBlock_3_0_2_0181_load_1),
        .p_read51(ap_sig_allocacmp_l_TBlock_3_0_3_0182_load_1),
        .p_read52(ap_sig_allocacmp_l_TBlock_3_1_0_0183_load_1),
        .p_read53(ap_sig_allocacmp_l_TBlock_3_1_1_0184_load_1),
        .p_read54(ap_sig_allocacmp_l_TBlock_3_1_2_0185_load_1),
        .p_read55(ap_sig_allocacmp_l_TBlock_3_1_3_0186_load_1),
        .p_read56(ap_sig_allocacmp_l_TBlock_3_2_0_0187_load_1),
        .p_read57(ap_sig_allocacmp_l_TBlock_3_2_1_0188_load_1),
        .p_read58(ap_sig_allocacmp_l_TBlock_3_2_2_0189_load_1),
        .p_read59(ap_sig_allocacmp_l_TBlock_3_2_3_0190_load_1),
        .p_read60(ap_sig_allocacmp_l_TBlock_3_3_0_0191_load_1),
        .p_read61(ap_sig_allocacmp_l_TBlock_3_3_1_0192_load_1),
        .p_read62(ap_sig_allocacmp_l_TBlock_3_3_2_0193_load_1),
        .p_read63(ap_sig_allocacmp_l_TBlock_3_3_3_0194_load_1),
        .H_offset(trunc_ln69_reg_2962),
        .ap_return_0(grp_rpyxyzToH_double_s_fu_984_ap_return_0),
        .ap_return_1(grp_rpyxyzToH_double_s_fu_984_ap_return_1),
        .ap_return_2(grp_rpyxyzToH_double_s_fu_984_ap_return_2),
        .ap_return_3(grp_rpyxyzToH_double_s_fu_984_ap_return_3),
        .ap_return_4(grp_rpyxyzToH_double_s_fu_984_ap_return_4),
        .ap_return_5(grp_rpyxyzToH_double_s_fu_984_ap_return_5),
        .ap_return_6(grp_rpyxyzToH_double_s_fu_984_ap_return_6),
        .ap_return_7(grp_rpyxyzToH_double_s_fu_984_ap_return_7),
        .ap_return_8(grp_rpyxyzToH_double_s_fu_984_ap_return_8),
        .ap_return_9(grp_rpyxyzToH_double_s_fu_984_ap_return_9),
        .ap_return_10(grp_rpyxyzToH_double_s_fu_984_ap_return_10),
        .ap_return_11(grp_rpyxyzToH_double_s_fu_984_ap_return_11),
        .ap_return_12(grp_rpyxyzToH_double_s_fu_984_ap_return_12),
        .ap_return_13(grp_rpyxyzToH_double_s_fu_984_ap_return_13),
        .ap_return_14(grp_rpyxyzToH_double_s_fu_984_ap_return_14),
        .ap_return_15(grp_rpyxyzToH_double_s_fu_984_ap_return_15),
        .ap_return_16(grp_rpyxyzToH_double_s_fu_984_ap_return_16),
        .ap_return_17(grp_rpyxyzToH_double_s_fu_984_ap_return_17),
        .ap_return_18(grp_rpyxyzToH_double_s_fu_984_ap_return_18),
        .ap_return_19(grp_rpyxyzToH_double_s_fu_984_ap_return_19),
        .ap_return_20(grp_rpyxyzToH_double_s_fu_984_ap_return_20),
        .ap_return_21(grp_rpyxyzToH_double_s_fu_984_ap_return_21),
        .ap_return_22(grp_rpyxyzToH_double_s_fu_984_ap_return_22),
        .ap_return_23(grp_rpyxyzToH_double_s_fu_984_ap_return_23),
        .ap_return_24(grp_rpyxyzToH_double_s_fu_984_ap_return_24),
        .ap_return_25(grp_rpyxyzToH_double_s_fu_984_ap_return_25),
        .ap_return_26(grp_rpyxyzToH_double_s_fu_984_ap_return_26),
        .ap_return_27(grp_rpyxyzToH_double_s_fu_984_ap_return_27),
        .ap_return_28(grp_rpyxyzToH_double_s_fu_984_ap_return_28),
        .ap_return_29(grp_rpyxyzToH_double_s_fu_984_ap_return_29),
        .ap_return_30(grp_rpyxyzToH_double_s_fu_984_ap_return_30),
        .ap_return_31(grp_rpyxyzToH_double_s_fu_984_ap_return_31),
        .ap_return_32(grp_rpyxyzToH_double_s_fu_984_ap_return_32),
        .ap_return_33(grp_rpyxyzToH_double_s_fu_984_ap_return_33),
        .ap_return_34(grp_rpyxyzToH_double_s_fu_984_ap_return_34),
        .ap_return_35(grp_rpyxyzToH_double_s_fu_984_ap_return_35),
        .ap_return_36(grp_rpyxyzToH_double_s_fu_984_ap_return_36),
        .ap_return_37(grp_rpyxyzToH_double_s_fu_984_ap_return_37),
        .ap_return_38(grp_rpyxyzToH_double_s_fu_984_ap_return_38),
        .ap_return_39(grp_rpyxyzToH_double_s_fu_984_ap_return_39),
        .ap_return_40(grp_rpyxyzToH_double_s_fu_984_ap_return_40),
        .ap_return_41(grp_rpyxyzToH_double_s_fu_984_ap_return_41),
        .ap_return_42(grp_rpyxyzToH_double_s_fu_984_ap_return_42),
        .ap_return_43(grp_rpyxyzToH_double_s_fu_984_ap_return_43),
        .ap_return_44(grp_rpyxyzToH_double_s_fu_984_ap_return_44),
        .ap_return_45(grp_rpyxyzToH_double_s_fu_984_ap_return_45),
        .ap_return_46(grp_rpyxyzToH_double_s_fu_984_ap_return_46),
        .ap_return_47(grp_rpyxyzToH_double_s_fu_984_ap_return_47),
        .ap_return_48(grp_rpyxyzToH_double_s_fu_984_ap_return_48),
        .ap_return_49(grp_rpyxyzToH_double_s_fu_984_ap_return_49),
        .ap_return_50(grp_rpyxyzToH_double_s_fu_984_ap_return_50),
        .ap_return_51(grp_rpyxyzToH_double_s_fu_984_ap_return_51),
        .ap_return_52(grp_rpyxyzToH_double_s_fu_984_ap_return_52),
        .ap_return_53(grp_rpyxyzToH_double_s_fu_984_ap_return_53),
        .ap_return_54(grp_rpyxyzToH_double_s_fu_984_ap_return_54),
        .ap_return_55(grp_rpyxyzToH_double_s_fu_984_ap_return_55),
        .ap_return_56(grp_rpyxyzToH_double_s_fu_984_ap_return_56),
        .ap_return_57(grp_rpyxyzToH_double_s_fu_984_ap_return_57),
        .ap_return_58(grp_rpyxyzToH_double_s_fu_984_ap_return_58),
        .ap_return_59(grp_rpyxyzToH_double_s_fu_984_ap_return_59),
        .ap_return_60(grp_rpyxyzToH_double_s_fu_984_ap_return_60),
        .ap_return_61(grp_rpyxyzToH_double_s_fu_984_ap_return_61),
        .ap_return_62(grp_rpyxyzToH_double_s_fu_984_ap_return_62),
        .ap_return_63(grp_rpyxyzToH_double_s_fu_984_ap_return_63)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U706 (
        .din0(64'd0),
        .din1(64'd4590068740216009523),
        .din2(64'd4583439441564520153),
        .din3(64'd4588087156379966505),
        .din4(trunc_ln69_fu_1076_p1),
        .dout(tmp_fu_1080_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U707 (
        .din0(64'd0),
        .din1(64'd0),
        .din2(64'd13801443187663470330),
        .din3(64'd0),
        .din4(trunc_ln69_fu_1076_p1),
        .dout(tmp_s_fu_1094_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U708 (
        .din0(64'd4591149604126578442),
        .din1(64'd0),
        .din2(64'd0),
        .din3(64'd4576918229304087675),
        .din4(trunc_ln69_fu_1076_p1),
        .dout(tmp_270_fu_1108_p6)
    );

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage1),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage1)) begin
                ap_enable_reg_pp0_iter0_reg <= 1'b0;
            end else if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b1 == ap_CS_fsm_pp0_stage77) & (1'b0 == ap_block_pp0_stage77_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln69_fu_1064_p2 == 1'd0))) begin
                i_1_fu_276 <= add_ln69_fu_1070_p2;
            end else if ((ap_loop_init == 1'b1)) begin
                i_1_fu_276 <= 3'd0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            icmp_ln69_reg_2958 <= icmp_ln69_fu_1064_p2;
            tmp_270_reg_2977 <= tmp_270_fu_1108_p6;
            tmp_reg_2967 <= tmp_fu_1080_p6;
            tmp_s_reg_2972 <= tmp_s_fu_1094_p6;
            trunc_ln69_reg_2962 <= trunc_ln69_fu_1076_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_0_0_0131_fu_280 <= grp_rpyxyzToH_double_s_fu_984_ap_return_0;
            l_TBlock_0_0_1_0132_fu_284 <= grp_rpyxyzToH_double_s_fu_984_ap_return_1;
            l_TBlock_0_0_2_0133_fu_288 <= grp_rpyxyzToH_double_s_fu_984_ap_return_2;
            l_TBlock_0_0_3_0134_fu_292 <= grp_rpyxyzToH_double_s_fu_984_ap_return_3;
            l_TBlock_0_1_0_0135_fu_296 <= grp_rpyxyzToH_double_s_fu_984_ap_return_4;
            l_TBlock_0_1_1_0136_fu_300 <= grp_rpyxyzToH_double_s_fu_984_ap_return_5;
            l_TBlock_0_1_2_0137_fu_304 <= grp_rpyxyzToH_double_s_fu_984_ap_return_6;
            l_TBlock_0_1_3_0138_fu_308 <= grp_rpyxyzToH_double_s_fu_984_ap_return_7;
            l_TBlock_0_2_0_0139_fu_312 <= grp_rpyxyzToH_double_s_fu_984_ap_return_8;
            l_TBlock_0_2_1_0140_fu_316 <= grp_rpyxyzToH_double_s_fu_984_ap_return_9;
            l_TBlock_0_2_2_0141_fu_320 <= grp_rpyxyzToH_double_s_fu_984_ap_return_10;
            l_TBlock_0_2_3_0142_fu_324 <= grp_rpyxyzToH_double_s_fu_984_ap_return_11;
            l_TBlock_0_3_0_0143_fu_328 <= grp_rpyxyzToH_double_s_fu_984_ap_return_12;
            l_TBlock_0_3_1_0144_fu_332 <= grp_rpyxyzToH_double_s_fu_984_ap_return_13;
            l_TBlock_0_3_2_0145_fu_336 <= grp_rpyxyzToH_double_s_fu_984_ap_return_14;
            l_TBlock_0_3_3_0146_fu_340 <= grp_rpyxyzToH_double_s_fu_984_ap_return_15;
            l_TBlock_1_0_0_0147_fu_344 <= grp_rpyxyzToH_double_s_fu_984_ap_return_16;
            l_TBlock_1_0_1_0148_fu_348 <= grp_rpyxyzToH_double_s_fu_984_ap_return_17;
            l_TBlock_1_0_2_0149_fu_352 <= grp_rpyxyzToH_double_s_fu_984_ap_return_18;
            l_TBlock_1_0_3_0150_fu_356 <= grp_rpyxyzToH_double_s_fu_984_ap_return_19;
            l_TBlock_1_1_0_0151_fu_360 <= grp_rpyxyzToH_double_s_fu_984_ap_return_20;
            l_TBlock_1_1_1_0152_fu_364 <= grp_rpyxyzToH_double_s_fu_984_ap_return_21;
            l_TBlock_1_1_2_0153_fu_368 <= grp_rpyxyzToH_double_s_fu_984_ap_return_22;
            l_TBlock_1_1_3_0154_fu_372 <= grp_rpyxyzToH_double_s_fu_984_ap_return_23;
            l_TBlock_1_2_0_0155_fu_376 <= grp_rpyxyzToH_double_s_fu_984_ap_return_24;
            l_TBlock_1_2_1_0156_fu_380 <= grp_rpyxyzToH_double_s_fu_984_ap_return_25;
            l_TBlock_1_2_2_0157_fu_384 <= grp_rpyxyzToH_double_s_fu_984_ap_return_26;
            l_TBlock_1_2_3_0158_fu_388 <= grp_rpyxyzToH_double_s_fu_984_ap_return_27;
            l_TBlock_1_3_0_0159_fu_392 <= grp_rpyxyzToH_double_s_fu_984_ap_return_28;
            l_TBlock_1_3_1_0160_fu_396 <= grp_rpyxyzToH_double_s_fu_984_ap_return_29;
            l_TBlock_1_3_2_0161_fu_400 <= grp_rpyxyzToH_double_s_fu_984_ap_return_30;
            l_TBlock_1_3_3_0162_fu_404 <= grp_rpyxyzToH_double_s_fu_984_ap_return_31;
            l_TBlock_2_0_0_0163_fu_408 <= grp_rpyxyzToH_double_s_fu_984_ap_return_32;
            l_TBlock_2_0_1_0164_fu_412 <= grp_rpyxyzToH_double_s_fu_984_ap_return_33;
            l_TBlock_2_0_2_0165_fu_416 <= grp_rpyxyzToH_double_s_fu_984_ap_return_34;
            l_TBlock_2_0_3_0166_fu_420 <= grp_rpyxyzToH_double_s_fu_984_ap_return_35;
            l_TBlock_2_1_0_0167_fu_424 <= grp_rpyxyzToH_double_s_fu_984_ap_return_36;
            l_TBlock_2_1_1_0168_fu_428 <= grp_rpyxyzToH_double_s_fu_984_ap_return_37;
            l_TBlock_2_1_2_0169_fu_432 <= grp_rpyxyzToH_double_s_fu_984_ap_return_38;
            l_TBlock_2_1_3_0170_fu_436 <= grp_rpyxyzToH_double_s_fu_984_ap_return_39;
            l_TBlock_2_2_0_0171_fu_440 <= grp_rpyxyzToH_double_s_fu_984_ap_return_40;
            l_TBlock_2_2_1_0172_fu_444 <= grp_rpyxyzToH_double_s_fu_984_ap_return_41;
            l_TBlock_2_2_2_0173_fu_448 <= grp_rpyxyzToH_double_s_fu_984_ap_return_42;
            l_TBlock_2_2_3_0174_fu_452 <= grp_rpyxyzToH_double_s_fu_984_ap_return_43;
            l_TBlock_2_3_0_0175_fu_456 <= grp_rpyxyzToH_double_s_fu_984_ap_return_44;
            l_TBlock_2_3_1_0176_fu_460 <= grp_rpyxyzToH_double_s_fu_984_ap_return_45;
            l_TBlock_2_3_2_0177_fu_464 <= grp_rpyxyzToH_double_s_fu_984_ap_return_46;
            l_TBlock_2_3_3_0178_fu_468 <= grp_rpyxyzToH_double_s_fu_984_ap_return_47;
            l_TBlock_3_0_0_0179_fu_472 <= grp_rpyxyzToH_double_s_fu_984_ap_return_48;
            l_TBlock_3_0_1_0180_fu_476 <= grp_rpyxyzToH_double_s_fu_984_ap_return_49;
            l_TBlock_3_0_2_0181_fu_480 <= grp_rpyxyzToH_double_s_fu_984_ap_return_50;
            l_TBlock_3_0_3_0182_fu_484 <= grp_rpyxyzToH_double_s_fu_984_ap_return_51;
            l_TBlock_3_1_0_0183_fu_488 <= grp_rpyxyzToH_double_s_fu_984_ap_return_52;
            l_TBlock_3_1_1_0184_fu_492 <= grp_rpyxyzToH_double_s_fu_984_ap_return_53;
            l_TBlock_3_1_2_0185_fu_496 <= grp_rpyxyzToH_double_s_fu_984_ap_return_54;
            l_TBlock_3_1_3_0186_fu_500 <= grp_rpyxyzToH_double_s_fu_984_ap_return_55;
            l_TBlock_3_2_0_0187_fu_504 <= grp_rpyxyzToH_double_s_fu_984_ap_return_56;
            l_TBlock_3_2_1_0188_fu_508 <= grp_rpyxyzToH_double_s_fu_984_ap_return_57;
            l_TBlock_3_2_2_0189_fu_512 <= grp_rpyxyzToH_double_s_fu_984_ap_return_58;
            l_TBlock_3_2_3_0190_fu_516 <= grp_rpyxyzToH_double_s_fu_984_ap_return_59;
            l_TBlock_3_3_0_0191_fu_520 <= grp_rpyxyzToH_double_s_fu_984_ap_return_60;
            l_TBlock_3_3_1_0192_fu_524 <= grp_rpyxyzToH_double_s_fu_984_ap_return_61;
            l_TBlock_3_3_2_0193_fu_528 <= grp_rpyxyzToH_double_s_fu_984_ap_return_62;
            l_TBlock_3_3_3_0194_fu_532 <= grp_rpyxyzToH_double_s_fu_984_ap_return_63;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_condition_exit_pp0_iter0_stage1 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_idle_pp0 == 1'b1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b0)) begin
            ap_idle_pp0_1to1 = 1'b1;
        end else begin
            ap_idle_pp0_1to1 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage77) & (1'b0 == ap_block_pp0_stage77_subdone))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ap_sig_allocacmp_i = 3'd0;
        end else begin
            ap_sig_allocacmp_i = i_1_fu_276;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_0_0_0131_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_0;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_0_0_0131_load_1 = l_TBlock_0_0_0_0131_fu_280;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_0_1_0132_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_1;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_0_1_0132_load_1 = l_TBlock_0_0_1_0132_fu_284;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_0_2_0133_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_2;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_0_2_0133_load_1 = l_TBlock_0_0_2_0133_fu_288;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_0_3_0134_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_3;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_0_3_0134_load_1 = l_TBlock_0_0_3_0134_fu_292;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_1_0_0135_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_4;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_1_0_0135_load_1 = l_TBlock_0_1_0_0135_fu_296;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_1_1_0136_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_5;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_1_1_0136_load_1 = l_TBlock_0_1_1_0136_fu_300;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_1_2_0137_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_6;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_1_2_0137_load_1 = l_TBlock_0_1_2_0137_fu_304;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_1_3_0138_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_7;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_1_3_0138_load_1 = l_TBlock_0_1_3_0138_fu_308;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_2_0_0139_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_8;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_2_0_0139_load_1 = l_TBlock_0_2_0_0139_fu_312;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_2_1_0140_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_9;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_2_1_0140_load_1 = l_TBlock_0_2_1_0140_fu_316;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_2_2_0141_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_10;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_2_2_0141_load_1 = l_TBlock_0_2_2_0141_fu_320;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_2_3_0142_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_11;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_2_3_0142_load_1 = l_TBlock_0_2_3_0142_fu_324;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_3_0_0143_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_12;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_3_0_0143_load_1 = l_TBlock_0_3_0_0143_fu_328;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_3_1_0144_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_13;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_3_1_0144_load_1 = l_TBlock_0_3_1_0144_fu_332;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_3_2_0145_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_14;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_3_2_0145_load_1 = l_TBlock_0_3_2_0145_fu_336;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_0_3_3_0146_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_15;
        end else begin
            ap_sig_allocacmp_l_TBlock_0_3_3_0146_load_1 = l_TBlock_0_3_3_0146_fu_340;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_0_0_0147_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_16;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_0_0_0147_load_1 = l_TBlock_1_0_0_0147_fu_344;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_0_1_0148_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_17;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_0_1_0148_load_1 = l_TBlock_1_0_1_0148_fu_348;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_0_2_0149_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_18;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_0_2_0149_load_1 = l_TBlock_1_0_2_0149_fu_352;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_0_3_0150_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_19;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_0_3_0150_load_1 = l_TBlock_1_0_3_0150_fu_356;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_1_0_0151_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_20;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_1_0_0151_load_1 = l_TBlock_1_1_0_0151_fu_360;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_1_1_0152_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_21;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_1_1_0152_load_1 = l_TBlock_1_1_1_0152_fu_364;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_1_2_0153_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_22;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_1_2_0153_load_1 = l_TBlock_1_1_2_0153_fu_368;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_1_3_0154_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_23;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_1_3_0154_load_1 = l_TBlock_1_1_3_0154_fu_372;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_2_0_0155_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_24;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_2_0_0155_load_1 = l_TBlock_1_2_0_0155_fu_376;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_2_1_0156_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_25;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_2_1_0156_load_1 = l_TBlock_1_2_1_0156_fu_380;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_2_2_0157_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_26;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_2_2_0157_load_1 = l_TBlock_1_2_2_0157_fu_384;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_2_3_0158_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_27;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_2_3_0158_load_1 = l_TBlock_1_2_3_0158_fu_388;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_3_0_0159_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_28;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_3_0_0159_load_1 = l_TBlock_1_3_0_0159_fu_392;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_3_1_0160_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_29;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_3_1_0160_load_1 = l_TBlock_1_3_1_0160_fu_396;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_3_2_0161_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_30;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_3_2_0161_load_1 = l_TBlock_1_3_2_0161_fu_400;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_1_3_3_0162_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_31;
        end else begin
            ap_sig_allocacmp_l_TBlock_1_3_3_0162_load_1 = l_TBlock_1_3_3_0162_fu_404;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_0_0_0163_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_32;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_0_0_0163_load_1 = l_TBlock_2_0_0_0163_fu_408;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_0_1_0164_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_33;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_0_1_0164_load_1 = l_TBlock_2_0_1_0164_fu_412;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_0_2_0165_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_34;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_0_2_0165_load_1 = l_TBlock_2_0_2_0165_fu_416;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_0_3_0166_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_35;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_0_3_0166_load_1 = l_TBlock_2_0_3_0166_fu_420;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_1_0_0167_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_36;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_1_0_0167_load_1 = l_TBlock_2_1_0_0167_fu_424;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_1_1_0168_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_37;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_1_1_0168_load_1 = l_TBlock_2_1_1_0168_fu_428;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_1_2_0169_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_38;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_1_2_0169_load_1 = l_TBlock_2_1_2_0169_fu_432;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_1_3_0170_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_39;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_1_3_0170_load_1 = l_TBlock_2_1_3_0170_fu_436;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_2_0_0171_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_40;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_2_0_0171_load_1 = l_TBlock_2_2_0_0171_fu_440;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_2_1_0172_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_41;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_2_1_0172_load_1 = l_TBlock_2_2_1_0172_fu_444;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_2_2_0173_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_42;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_2_2_0173_load_1 = l_TBlock_2_2_2_0173_fu_448;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_2_3_0174_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_43;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_2_3_0174_load_1 = l_TBlock_2_2_3_0174_fu_452;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_3_0_0175_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_44;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_3_0_0175_load_1 = l_TBlock_2_3_0_0175_fu_456;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_3_1_0176_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_45;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_3_1_0176_load_1 = l_TBlock_2_3_1_0176_fu_460;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_3_2_0177_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_46;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_3_2_0177_load_1 = l_TBlock_2_3_2_0177_fu_464;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_2_3_3_0178_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_47;
        end else begin
            ap_sig_allocacmp_l_TBlock_2_3_3_0178_load_1 = l_TBlock_2_3_3_0178_fu_468;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_0_0_0179_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_48;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_0_0_0179_load_1 = l_TBlock_3_0_0_0179_fu_472;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_0_1_0180_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_49;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_0_1_0180_load_1 = l_TBlock_3_0_1_0180_fu_476;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_0_2_0181_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_50;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_0_2_0181_load_1 = l_TBlock_3_0_2_0181_fu_480;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_0_3_0182_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_51;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_0_3_0182_load_1 = l_TBlock_3_0_3_0182_fu_484;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_1_0_0183_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_52;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_1_0_0183_load_1 = l_TBlock_3_1_0_0183_fu_488;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_1_1_0184_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_53;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_1_1_0184_load_1 = l_TBlock_3_1_1_0184_fu_492;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_1_2_0185_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_54;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_1_2_0185_load_1 = l_TBlock_3_1_2_0185_fu_496;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_1_3_0186_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_55;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_1_3_0186_load_1 = l_TBlock_3_1_3_0186_fu_500;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_2_0_0187_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_56;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_2_0_0187_load_1 = l_TBlock_3_2_0_0187_fu_504;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_2_1_0188_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_57;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_2_1_0188_load_1 = l_TBlock_3_2_1_0188_fu_508;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_2_2_0189_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_58;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_2_2_0189_load_1 = l_TBlock_3_2_2_0189_fu_512;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_2_3_0190_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_59;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_2_3_0190_load_1 = l_TBlock_3_2_3_0190_fu_516;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_3_0_0191_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_60;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_3_0_0191_load_1 = l_TBlock_3_3_0_0191_fu_520;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_3_1_0192_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_61;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_3_1_0192_load_1 = l_TBlock_3_3_1_0192_fu_524;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_3_2_0193_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_62;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_3_2_0193_load_1 = l_TBlock_3_3_2_0193_fu_528;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ap_sig_allocacmp_l_TBlock_3_3_3_0194_load_1 = grp_rpyxyzToH_double_s_fu_984_ap_return_63;
        end else begin
            ap_sig_allocacmp_l_TBlock_3_3_3_0194_load_1 = l_TBlock_3_3_3_0194_fu_532;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_0_0_0131_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_0_0_0131_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_0_1_0132_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_0_1_0132_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_0_2_0133_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_0_2_0133_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_0_3_0134_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_0_3_0134_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_1_0_0135_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_1_0_0135_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_1_1_0136_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_1_1_0136_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_1_2_0137_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_1_2_0137_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_1_3_0138_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_1_3_0138_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_2_0_0139_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_2_0_0139_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_2_1_0140_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_2_1_0140_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_2_2_0141_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_2_2_0141_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_2_3_0142_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_2_3_0142_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_3_0_0143_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_3_0_0143_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_3_1_0144_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_3_1_0144_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_3_2_0145_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_3_2_0145_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_0_3_3_0146_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_0_3_3_0146_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_0_0_0147_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_0_0_0147_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_0_1_0148_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_0_1_0148_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_0_2_0149_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_0_2_0149_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_0_3_0150_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_0_3_0150_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_1_0_0151_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_1_0_0151_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_1_1_0152_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_1_1_0152_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_1_2_0153_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_1_2_0153_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_1_3_0154_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_1_3_0154_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_2_0_0155_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_2_0_0155_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_2_1_0156_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_2_1_0156_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_2_2_0157_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_2_2_0157_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_2_3_0158_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_2_3_0158_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_3_0_0159_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_3_0_0159_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_3_1_0160_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_3_1_0160_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_3_2_0161_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_3_2_0161_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_1_3_3_0162_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_1_3_3_0162_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_0_0_0163_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_0_0_0163_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_0_1_0164_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_0_1_0164_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_0_2_0165_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_0_2_0165_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_0_3_0166_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_0_3_0166_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_1_0_0167_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_1_0_0167_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_1_1_0168_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_1_1_0168_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_1_2_0169_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_1_2_0169_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_1_3_0170_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_1_3_0170_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_2_0_0171_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_2_0_0171_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_2_1_0172_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_2_1_0172_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_2_2_0173_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_2_2_0173_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_2_3_0174_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_2_3_0174_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_3_0_0175_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_3_0_0175_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_3_1_0176_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_3_1_0176_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_3_2_0177_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_3_2_0177_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_2_3_3_0178_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_2_3_3_0178_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_0_0_0179_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_0_0_0179_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_0_1_0180_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_0_1_0180_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_0_2_0181_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_0_2_0181_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_0_3_0182_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_0_3_0182_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_1_0_0183_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_1_0_0183_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_1_1_0184_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_1_1_0184_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_1_2_0185_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_1_2_0185_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_1_3_0186_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_1_3_0186_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_2_0_0187_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_2_0_0187_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_2_1_0188_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_2_1_0188_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_2_2_0189_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_2_2_0189_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_2_3_0190_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_2_3_0190_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_3_0_0191_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_3_0_0191_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_3_1_0192_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_3_1_0192_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_3_2_0193_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_3_2_0193_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln69_reg_2958 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
            l_TBlock_3_3_3_0194_out_ap_vld = 1'b1;
        end else begin
            l_TBlock_3_3_3_0194_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_0_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_0_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_0_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_0_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_0_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_1_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_1_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_1_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_1_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_1_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_2_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_2_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_2_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_2_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_2_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_3_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_3_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_3_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_0_3_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_0_3_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_0_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_0_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_0_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_0_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_0_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_1_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_1_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_1_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_1_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_1_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_2_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_2_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_2_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_2_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_2_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_3_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_3_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_3_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_1_3_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_1_3_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_0_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_0_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_0_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_0_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_0_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_1_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_1_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_1_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_1_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_1_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_2_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_2_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_2_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_2_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_2_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd0) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_3_0_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_0_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd1) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_3_1_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_1_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd2) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_3_2_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_2_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (trunc_ln69_fu_1076_p1 == 2'd3) & (icmp_ln69_fu_1064_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            l_TColl_2_3_3_constprop_ap_vld = 1'b1;
        end else begin
            l_TColl_2_3_3_constprop_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to1 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b1 == ap_condition_exit_pp0_iter0_stage1)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if ((1'b0 == ap_block_pp0_stage9_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            ap_ST_fsm_pp0_stage14: begin
                if ((1'b0 == ap_block_pp0_stage14_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage14;
                end
            end
            ap_ST_fsm_pp0_stage15: begin
                if ((1'b0 == ap_block_pp0_stage15_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage15;
                end
            end
            ap_ST_fsm_pp0_stage16: begin
                if ((1'b0 == ap_block_pp0_stage16_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage16;
                end
            end
            ap_ST_fsm_pp0_stage17: begin
                if ((1'b0 == ap_block_pp0_stage17_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage17;
                end
            end
            ap_ST_fsm_pp0_stage18: begin
                if ((1'b0 == ap_block_pp0_stage18_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage18;
                end
            end
            ap_ST_fsm_pp0_stage19: begin
                if ((1'b0 == ap_block_pp0_stage19_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage19;
                end
            end
            ap_ST_fsm_pp0_stage20: begin
                if ((1'b0 == ap_block_pp0_stage20_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage20;
                end
            end
            ap_ST_fsm_pp0_stage21: begin
                if ((1'b0 == ap_block_pp0_stage21_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage21;
                end
            end
            ap_ST_fsm_pp0_stage22: begin
                if ((1'b0 == ap_block_pp0_stage22_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage22;
                end
            end
            ap_ST_fsm_pp0_stage23: begin
                if ((1'b0 == ap_block_pp0_stage23_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage23;
                end
            end
            ap_ST_fsm_pp0_stage24: begin
                if ((1'b0 == ap_block_pp0_stage24_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage24;
                end
            end
            ap_ST_fsm_pp0_stage25: begin
                if ((1'b0 == ap_block_pp0_stage25_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage25;
                end
            end
            ap_ST_fsm_pp0_stage26: begin
                if ((1'b0 == ap_block_pp0_stage26_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage26;
                end
            end
            ap_ST_fsm_pp0_stage27: begin
                if ((1'b0 == ap_block_pp0_stage27_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage27;
                end
            end
            ap_ST_fsm_pp0_stage28: begin
                if ((1'b0 == ap_block_pp0_stage28_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage28;
                end
            end
            ap_ST_fsm_pp0_stage29: begin
                if ((1'b0 == ap_block_pp0_stage29_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage29;
                end
            end
            ap_ST_fsm_pp0_stage30: begin
                if ((1'b0 == ap_block_pp0_stage30_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage30;
                end
            end
            ap_ST_fsm_pp0_stage31: begin
                if ((1'b0 == ap_block_pp0_stage31_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage31;
                end
            end
            ap_ST_fsm_pp0_stage32: begin
                if ((1'b0 == ap_block_pp0_stage32_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage32;
                end
            end
            ap_ST_fsm_pp0_stage33: begin
                if ((1'b0 == ap_block_pp0_stage33_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage33;
                end
            end
            ap_ST_fsm_pp0_stage34: begin
                if ((1'b0 == ap_block_pp0_stage34_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage34;
                end
            end
            ap_ST_fsm_pp0_stage35: begin
                if ((1'b0 == ap_block_pp0_stage35_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage35;
                end
            end
            ap_ST_fsm_pp0_stage36: begin
                if ((1'b0 == ap_block_pp0_stage36_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage36;
                end
            end
            ap_ST_fsm_pp0_stage37: begin
                if ((1'b0 == ap_block_pp0_stage37_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage37;
                end
            end
            ap_ST_fsm_pp0_stage38: begin
                if ((1'b0 == ap_block_pp0_stage38_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage38;
                end
            end
            ap_ST_fsm_pp0_stage39: begin
                if ((1'b0 == ap_block_pp0_stage39_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage39;
                end
            end
            ap_ST_fsm_pp0_stage40: begin
                if ((1'b0 == ap_block_pp0_stage40_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage40;
                end
            end
            ap_ST_fsm_pp0_stage41: begin
                if ((1'b0 == ap_block_pp0_stage41_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage41;
                end
            end
            ap_ST_fsm_pp0_stage42: begin
                if ((1'b0 == ap_block_pp0_stage42_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage42;
                end
            end
            ap_ST_fsm_pp0_stage43: begin
                if ((1'b0 == ap_block_pp0_stage43_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage43;
                end
            end
            ap_ST_fsm_pp0_stage44: begin
                if ((1'b0 == ap_block_pp0_stage44_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage44;
                end
            end
            ap_ST_fsm_pp0_stage45: begin
                if ((1'b0 == ap_block_pp0_stage45_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage45;
                end
            end
            ap_ST_fsm_pp0_stage46: begin
                if ((1'b0 == ap_block_pp0_stage46_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage46;
                end
            end
            ap_ST_fsm_pp0_stage47: begin
                if ((1'b0 == ap_block_pp0_stage47_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage47;
                end
            end
            ap_ST_fsm_pp0_stage48: begin
                if ((1'b0 == ap_block_pp0_stage48_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage48;
                end
            end
            ap_ST_fsm_pp0_stage49: begin
                if ((1'b0 == ap_block_pp0_stage49_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage49;
                end
            end
            ap_ST_fsm_pp0_stage50: begin
                if ((1'b0 == ap_block_pp0_stage50_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage50;
                end
            end
            ap_ST_fsm_pp0_stage51: begin
                if ((1'b0 == ap_block_pp0_stage51_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage51;
                end
            end
            ap_ST_fsm_pp0_stage52: begin
                if ((1'b0 == ap_block_pp0_stage52_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage52;
                end
            end
            ap_ST_fsm_pp0_stage53: begin
                if ((1'b0 == ap_block_pp0_stage53_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage53;
                end
            end
            ap_ST_fsm_pp0_stage54: begin
                if ((1'b0 == ap_block_pp0_stage54_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage54;
                end
            end
            ap_ST_fsm_pp0_stage55: begin
                if ((1'b0 == ap_block_pp0_stage55_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage55;
                end
            end
            ap_ST_fsm_pp0_stage56: begin
                if ((1'b0 == ap_block_pp0_stage56_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage56;
                end
            end
            ap_ST_fsm_pp0_stage57: begin
                if ((1'b0 == ap_block_pp0_stage57_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage57;
                end
            end
            ap_ST_fsm_pp0_stage58: begin
                if ((1'b0 == ap_block_pp0_stage58_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage58;
                end
            end
            ap_ST_fsm_pp0_stage59: begin
                if ((1'b0 == ap_block_pp0_stage59_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage59;
                end
            end
            ap_ST_fsm_pp0_stage60: begin
                if ((1'b0 == ap_block_pp0_stage60_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage60;
                end
            end
            ap_ST_fsm_pp0_stage61: begin
                if ((1'b0 == ap_block_pp0_stage61_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage61;
                end
            end
            ap_ST_fsm_pp0_stage62: begin
                if ((1'b0 == ap_block_pp0_stage62_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage62;
                end
            end
            ap_ST_fsm_pp0_stage63: begin
                if ((1'b0 == ap_block_pp0_stage63_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage63;
                end
            end
            ap_ST_fsm_pp0_stage64: begin
                if ((1'b0 == ap_block_pp0_stage64_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage64;
                end
            end
            ap_ST_fsm_pp0_stage65: begin
                if ((1'b0 == ap_block_pp0_stage65_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage65;
                end
            end
            ap_ST_fsm_pp0_stage66: begin
                if ((1'b0 == ap_block_pp0_stage66_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage66;
                end
            end
            ap_ST_fsm_pp0_stage67: begin
                if ((1'b0 == ap_block_pp0_stage67_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage67;
                end
            end
            ap_ST_fsm_pp0_stage68: begin
                if ((1'b0 == ap_block_pp0_stage68_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage69;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage68;
                end
            end
            ap_ST_fsm_pp0_stage69: begin
                if ((1'b0 == ap_block_pp0_stage69_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage70;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage69;
                end
            end
            ap_ST_fsm_pp0_stage70: begin
                if ((1'b0 == ap_block_pp0_stage70_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage71;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage70;
                end
            end
            ap_ST_fsm_pp0_stage71: begin
                if ((1'b0 == ap_block_pp0_stage71_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage72;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage71;
                end
            end
            ap_ST_fsm_pp0_stage72: begin
                if ((1'b0 == ap_block_pp0_stage72_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage73;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage72;
                end
            end
            ap_ST_fsm_pp0_stage73: begin
                if ((1'b0 == ap_block_pp0_stage73_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage74;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage73;
                end
            end
            ap_ST_fsm_pp0_stage74: begin
                if ((1'b0 == ap_block_pp0_stage74_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage75;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage74;
                end
            end
            ap_ST_fsm_pp0_stage75: begin
                if ((1'b0 == ap_block_pp0_stage75_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage76;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage75;
                end
            end
            ap_ST_fsm_pp0_stage76: begin
                if ((1'b0 == ap_block_pp0_stage76_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage77;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage76;
                end
            end
            ap_ST_fsm_pp0_stage77: begin
                if ((1'b0 == ap_block_pp0_stage77_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage77;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln69_fu_1070_p2 = (ap_sig_allocacmp_i + 3'd1);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage77 = ap_CS_fsm[32'd77];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage14_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage15_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage16_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage17_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage18_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage19_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage20_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage21_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage22_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage23_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage24_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage25_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage26_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage27_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage28_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage29_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage30_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage31_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage32_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage33_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage34_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage35_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage36_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage37_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage38_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage39_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage40_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage41_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage42_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage43_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage44_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage45_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage46_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage47_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage48_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage49_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage50_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage51_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage52_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage53_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage54_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage55_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage56_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage57_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage58_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage59_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage60_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage61_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage62_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage63_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage64_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage65_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage66_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage67_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage68_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage69_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage70_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage71_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage72_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage73_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage74_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage75_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage76_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage77_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage1;

    assign icmp_ln69_fu_1064_p2 = ((ap_sig_allocacmp_i == 3'd4) ? 1'b1 : 1'b0);

    assign l_TBlock_0_0_0_0131_out = l_TBlock_0_0_0_0131_fu_280;

    assign l_TBlock_0_0_1_0132_out = l_TBlock_0_0_1_0132_fu_284;

    assign l_TBlock_0_0_2_0133_out = l_TBlock_0_0_2_0133_fu_288;

    assign l_TBlock_0_0_3_0134_out = l_TBlock_0_0_3_0134_fu_292;

    assign l_TBlock_0_1_0_0135_out = l_TBlock_0_1_0_0135_fu_296;

    assign l_TBlock_0_1_1_0136_out = l_TBlock_0_1_1_0136_fu_300;

    assign l_TBlock_0_1_2_0137_out = l_TBlock_0_1_2_0137_fu_304;

    assign l_TBlock_0_1_3_0138_out = l_TBlock_0_1_3_0138_fu_308;

    assign l_TBlock_0_2_0_0139_out = l_TBlock_0_2_0_0139_fu_312;

    assign l_TBlock_0_2_1_0140_out = l_TBlock_0_2_1_0140_fu_316;

    assign l_TBlock_0_2_2_0141_out = l_TBlock_0_2_2_0141_fu_320;

    assign l_TBlock_0_2_3_0142_out = l_TBlock_0_2_3_0142_fu_324;

    assign l_TBlock_0_3_0_0143_out = l_TBlock_0_3_0_0143_fu_328;

    assign l_TBlock_0_3_1_0144_out = l_TBlock_0_3_1_0144_fu_332;

    assign l_TBlock_0_3_2_0145_out = l_TBlock_0_3_2_0145_fu_336;

    assign l_TBlock_0_3_3_0146_out = l_TBlock_0_3_3_0146_fu_340;

    assign l_TBlock_1_0_0_0147_out = l_TBlock_1_0_0_0147_fu_344;

    assign l_TBlock_1_0_1_0148_out = l_TBlock_1_0_1_0148_fu_348;

    assign l_TBlock_1_0_2_0149_out = l_TBlock_1_0_2_0149_fu_352;

    assign l_TBlock_1_0_3_0150_out = l_TBlock_1_0_3_0150_fu_356;

    assign l_TBlock_1_1_0_0151_out = l_TBlock_1_1_0_0151_fu_360;

    assign l_TBlock_1_1_1_0152_out = l_TBlock_1_1_1_0152_fu_364;

    assign l_TBlock_1_1_2_0153_out = l_TBlock_1_1_2_0153_fu_368;

    assign l_TBlock_1_1_3_0154_out = l_TBlock_1_1_3_0154_fu_372;

    assign l_TBlock_1_2_0_0155_out = l_TBlock_1_2_0_0155_fu_376;

    assign l_TBlock_1_2_1_0156_out = l_TBlock_1_2_1_0156_fu_380;

    assign l_TBlock_1_2_2_0157_out = l_TBlock_1_2_2_0157_fu_384;

    assign l_TBlock_1_2_3_0158_out = l_TBlock_1_2_3_0158_fu_388;

    assign l_TBlock_1_3_0_0159_out = l_TBlock_1_3_0_0159_fu_392;

    assign l_TBlock_1_3_1_0160_out = l_TBlock_1_3_1_0160_fu_396;

    assign l_TBlock_1_3_2_0161_out = l_TBlock_1_3_2_0161_fu_400;

    assign l_TBlock_1_3_3_0162_out = l_TBlock_1_3_3_0162_fu_404;

    assign l_TBlock_2_0_0_0163_out = l_TBlock_2_0_0_0163_fu_408;

    assign l_TBlock_2_0_1_0164_out = l_TBlock_2_0_1_0164_fu_412;

    assign l_TBlock_2_0_2_0165_out = l_TBlock_2_0_2_0165_fu_416;

    assign l_TBlock_2_0_3_0166_out = l_TBlock_2_0_3_0166_fu_420;

    assign l_TBlock_2_1_0_0167_out = l_TBlock_2_1_0_0167_fu_424;

    assign l_TBlock_2_1_1_0168_out = l_TBlock_2_1_1_0168_fu_428;

    assign l_TBlock_2_1_2_0169_out = l_TBlock_2_1_2_0169_fu_432;

    assign l_TBlock_2_1_3_0170_out = l_TBlock_2_1_3_0170_fu_436;

    assign l_TBlock_2_2_0_0171_out = l_TBlock_2_2_0_0171_fu_440;

    assign l_TBlock_2_2_1_0172_out = l_TBlock_2_2_1_0172_fu_444;

    assign l_TBlock_2_2_2_0173_out = l_TBlock_2_2_2_0173_fu_448;

    assign l_TBlock_2_2_3_0174_out = l_TBlock_2_2_3_0174_fu_452;

    assign l_TBlock_2_3_0_0175_out = l_TBlock_2_3_0_0175_fu_456;

    assign l_TBlock_2_3_1_0176_out = l_TBlock_2_3_1_0176_fu_460;

    assign l_TBlock_2_3_2_0177_out = l_TBlock_2_3_2_0177_fu_464;

    assign l_TBlock_2_3_3_0178_out = l_TBlock_2_3_3_0178_fu_468;

    assign l_TBlock_3_0_0_0179_out = l_TBlock_3_0_0_0179_fu_472;

    assign l_TBlock_3_0_1_0180_out = l_TBlock_3_0_1_0180_fu_476;

    assign l_TBlock_3_0_2_0181_out = l_TBlock_3_0_2_0181_fu_480;

    assign l_TBlock_3_0_3_0182_out = l_TBlock_3_0_3_0182_fu_484;

    assign l_TBlock_3_1_0_0183_out = l_TBlock_3_1_0_0183_fu_488;

    assign l_TBlock_3_1_1_0184_out = l_TBlock_3_1_1_0184_fu_492;

    assign l_TBlock_3_1_2_0185_out = l_TBlock_3_1_2_0185_fu_496;

    assign l_TBlock_3_1_3_0186_out = l_TBlock_3_1_3_0186_fu_500;

    assign l_TBlock_3_2_0_0187_out = l_TBlock_3_2_0_0187_fu_504;

    assign l_TBlock_3_2_1_0188_out = l_TBlock_3_2_1_0188_fu_508;

    assign l_TBlock_3_2_2_0189_out = l_TBlock_3_2_2_0189_fu_512;

    assign l_TBlock_3_2_3_0190_out = l_TBlock_3_2_3_0190_fu_516;

    assign l_TBlock_3_3_0_0191_out = l_TBlock_3_3_0_0191_fu_520;

    assign l_TBlock_3_3_1_0192_out = l_TBlock_3_3_1_0192_fu_524;

    assign l_TBlock_3_3_2_0193_out = l_TBlock_3_3_2_0193_fu_528;

    assign l_TBlock_3_3_3_0194_out = l_TBlock_3_3_3_0194_fu_532;

    assign l_TColl_0_0_0_constprop = 64'd4607182418800017408;

    assign l_TColl_0_0_1_constprop = 64'd4607182418800017408;

    assign l_TColl_0_0_2_constprop = 64'd4607182418800017408;

    assign l_TColl_0_0_3_constprop = 64'd4607182418800017408;

    assign l_TColl_0_1_0_constprop = 64'd0;

    assign l_TColl_0_1_1_constprop = 64'd0;

    assign l_TColl_0_1_2_constprop = 64'd0;

    assign l_TColl_0_1_3_constprop = 64'd0;

    assign l_TColl_0_2_0_constprop = 64'd0;

    assign l_TColl_0_2_1_constprop = 64'd0;

    assign l_TColl_0_2_2_constprop = 64'd0;

    assign l_TColl_0_2_3_constprop = 64'd0;

    assign l_TColl_0_3_0_constprop = 64'd0;

    assign l_TColl_0_3_1_constprop = 64'd0;

    assign l_TColl_0_3_2_constprop = 64'd0;

    assign l_TColl_0_3_3_constprop = 64'd0;

    assign l_TColl_1_0_0_constprop = 64'd0;

    assign l_TColl_1_0_1_constprop = 64'd0;

    assign l_TColl_1_0_2_constprop = 64'd0;

    assign l_TColl_1_0_3_constprop = 64'd0;

    assign l_TColl_1_1_0_constprop = 64'd4607182418800017408;

    assign l_TColl_1_1_1_constprop = 64'd4607182418800017408;

    assign l_TColl_1_1_2_constprop = 64'd4607182418800017408;

    assign l_TColl_1_1_3_constprop = 64'd4607182418800017408;

    assign l_TColl_1_2_0_constprop = 64'd0;

    assign l_TColl_1_2_1_constprop = 64'd0;

    assign l_TColl_1_2_2_constprop = 64'd0;

    assign l_TColl_1_2_3_constprop = 64'd0;

    assign l_TColl_1_3_0_constprop = 64'd0;

    assign l_TColl_1_3_1_constprop = 64'd0;

    assign l_TColl_1_3_2_constprop = 64'd0;

    assign l_TColl_1_3_3_constprop = 64'd0;

    assign l_TColl_2_0_0_constprop = 64'd0;

    assign l_TColl_2_0_1_constprop = 64'd0;

    assign l_TColl_2_0_2_constprop = 64'd0;

    assign l_TColl_2_0_3_constprop = 64'd0;

    assign l_TColl_2_1_0_constprop = 64'd0;

    assign l_TColl_2_1_1_constprop = 64'd0;

    assign l_TColl_2_1_2_constprop = 64'd0;

    assign l_TColl_2_1_3_constprop = 64'd0;

    assign l_TColl_2_2_0_constprop = 64'd4607182418800017408;

    assign l_TColl_2_2_1_constprop = 64'd4607182418800017408;

    assign l_TColl_2_2_2_constprop = 64'd4607182418800017408;

    assign l_TColl_2_2_3_constprop = 64'd4607182418800017408;

    assign l_TColl_2_3_0_constprop = 64'd0;

    assign l_TColl_2_3_1_constprop = 64'd0;

    assign l_TColl_2_3_2_constprop = 64'd0;

    assign l_TColl_2_3_3_constprop = 64'd0;

    assign trunc_ln69_fu_1076_p1 = ap_sig_allocacmp_i[1:0];

endmodule  //main_main_Pipeline_VITIS_LOOP_69_4
