/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_updateMotion_Pipeline_VITIS_LOOP_46_2 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    angle_assign_1_reload,
    angle_assign_3_out,
    angle_assign_3_out_ap_vld,
    grp_fu_323_p_din0,
    grp_fu_323_p_din1,
    grp_fu_323_p_opcode,
    grp_fu_323_p_dout0,
    grp_fu_323_p_ce,
    grp_fu_361_p_din0,
    grp_fu_361_p_din1,
    grp_fu_361_p_opcode,
    grp_fu_361_p_dout0,
    grp_fu_361_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 8'd1;
    parameter ap_ST_fsm_pp0_stage1 = 8'd2;
    parameter ap_ST_fsm_pp0_stage2 = 8'd4;
    parameter ap_ST_fsm_pp0_stage3 = 8'd8;
    parameter ap_ST_fsm_pp0_stage4 = 8'd16;
    parameter ap_ST_fsm_pp0_stage5 = 8'd32;
    parameter ap_ST_fsm_pp0_stage6 = 8'd64;
    parameter ap_ST_fsm_pp0_stage7 = 8'd128;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] angle_assign_1_reload;
    output [63:0] angle_assign_3_out;
    output angle_assign_3_out_ap_vld;
    output [63:0] grp_fu_323_p_din0;
    output [63:0] grp_fu_323_p_din1;
    output [0:0] grp_fu_323_p_opcode;
    input [63:0] grp_fu_323_p_dout0;
    output grp_fu_323_p_ce;
    output [63:0] grp_fu_361_p_din0;
    output [63:0] grp_fu_361_p_din1;
    output [4:0] grp_fu_361_p_opcode;
    input [0:0] grp_fu_361_p_dout0;
    output grp_fu_361_p_ce;

    reg ap_idle;
    reg angle_assign_3_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [7:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_subdone;
    wire   [0:0] and_ln46_fu_107_p2;
    reg    ap_condition_exit_pp0_iter0_stage2;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] angle_assign_3_load_reg_124;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire    ap_block_pp0_stage2_11001;
    reg   [63:0] angle_assign_4_reg_136;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage1_subdone;
    reg   [63:0] angle_assign_3_fu_36;
    reg   [63:0] ap_sig_allocacmp_angle_assign_3_load;
    wire    ap_block_pp0_stage1;
    wire    ap_loop_init;
    wire    ap_block_pp0_stage2_01001;
    wire    ap_block_pp0_stage0;
    wire    ap_block_pp0_stage2;
    wire   [63:0] bitcast_ln46_fu_72_p1;
    wire   [10:0] tmp_s_fu_75_p4;
    wire   [51:0] trunc_ln46_fu_85_p1;
    wire   [0:0] icmp_ln46_1_fu_95_p2;
    wire   [0:0] icmp_ln46_fu_89_p2;
    wire   [0:0] or_ln46_fu_101_p2;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage1_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg   [7:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to1;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 8'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 angle_assign_3_fu_36 = 64'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage2),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_condition_exit_pp0_iter0_stage2)) begin
                ap_enable_reg_pp0_iter0_reg <= 1'b0;
            end else if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                ap_enable_reg_pp0_iter1 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            angle_assign_3_fu_36 <= angle_assign_1_reload;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            angle_assign_3_fu_36 <= angle_assign_4_reg_136;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            angle_assign_3_load_reg_124 <= ap_sig_allocacmp_angle_assign_3_load;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            angle_assign_4_reg_136 <= grp_fu_323_p_dout0;
        end
    end

    always @(*) begin
        if (((1'd0 == and_ln46_fu_107_p2) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            angle_assign_3_out_ap_vld = 1'b1;
        end else begin
            angle_assign_3_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((1'd0 == and_ln46_fu_107_p2) & (1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_condition_exit_pp0_iter0_stage2 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage2 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter1 == 1'b0)) begin
            ap_idle_pp0_1to1 = 1'b1;
        end else begin
            ap_idle_pp0_1to1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage7_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_sig_allocacmp_angle_assign_3_load = angle_assign_4_reg_136;
        end else begin
            ap_sig_allocacmp_angle_assign_3_load = angle_assign_3_fu_36;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to1 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b1 == ap_condition_exit_pp0_iter0_stage2)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign and_ln46_fu_107_p2 = (or_ln46_fu_101_p2 & grp_fu_361_p_dout0);

    assign angle_assign_3_out = angle_assign_3_load_reg_124;

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage2;

    assign bitcast_ln46_fu_72_p1 = angle_assign_3_load_reg_124;

    assign grp_fu_323_p_ce = 1'b1;

    assign grp_fu_323_p_din0 = angle_assign_3_load_reg_124;

    assign grp_fu_323_p_din1 = 64'd4618760256180340048;

    assign grp_fu_323_p_opcode = 2'd0;

    assign grp_fu_361_p_ce = 1'b1;

    assign grp_fu_361_p_din0 = ap_sig_allocacmp_angle_assign_3_load;

    assign grp_fu_361_p_din1 = 64'd13837628693407745360;

    assign grp_fu_361_p_opcode = 5'd4;

    assign icmp_ln46_1_fu_95_p2 = ((trunc_ln46_fu_85_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln46_fu_89_p2 = ((tmp_s_fu_75_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign or_ln46_fu_101_p2 = (icmp_ln46_fu_89_p2 | icmp_ln46_1_fu_95_p2);

    assign tmp_s_fu_75_p4 = {{bitcast_ln46_fu_72_p1[62:52]}};

    assign trunc_ln46_fu_85_p1 = bitcast_ln46_fu_72_p1[51:0];

endmodule  //main_updateMotion_Pipeline_VITIS_LOOP_46_2
