/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_sin_or_cos_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    ap_ce,
    t_in,
    do_cos,
    ap_return
);

    parameter ap_ST_fsm_pp0_stage0 = 1'd1;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input ap_ce;
    input [63:0] t_in;
    input [0:0] do_cos;
    output [63:0] ap_return;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;

    (* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    wire    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_enable_reg_pp0_iter10;
    reg    ap_enable_reg_pp0_iter11;
    reg    ap_enable_reg_pp0_iter12;
    reg    ap_enable_reg_pp0_iter13;
    reg    ap_enable_reg_pp0_iter14;
    reg    ap_enable_reg_pp0_iter15;
    reg    ap_enable_reg_pp0_iter16;
    reg    ap_enable_reg_pp0_iter17;
    reg    ap_enable_reg_pp0_iter18;
    reg    ap_enable_reg_pp0_iter19;
    reg    ap_enable_reg_pp0_iter20;
    reg    ap_enable_reg_pp0_iter21;
    reg    ap_enable_reg_pp0_iter22;
    reg    ap_enable_reg_pp0_iter23;
    reg    ap_enable_reg_pp0_iter24;
    reg    ap_enable_reg_pp0_iter25;
    reg    ap_enable_reg_pp0_iter26;
    reg    ap_enable_reg_pp0_iter27;
    reg    ap_enable_reg_pp0_iter28;
    reg    ap_enable_reg_pp0_iter29;
    reg    ap_enable_reg_pp0_iter30;
    reg    ap_enable_reg_pp0_iter31;
    reg    ap_enable_reg_pp0_iter32;
    reg    ap_idle_pp0;
    reg    ap_block_pp0_stage0_subdone;
    wire   [3:0] ref_4oPi_table_256_address0;
    reg    ref_4oPi_table_256_ce0;
    wire   [255:0] ref_4oPi_table_256_q0;
    wire   [7:0] fourth_order_double_sin_cos_K0_address0;
    reg    fourth_order_double_sin_cos_K0_ce0;
    wire   [58:0] fourth_order_double_sin_cos_K0_q0;
    wire   [7:0] fourth_order_double_sin_cos_K1_address0;
    reg    fourth_order_double_sin_cos_K1_ce0;
    wire   [51:0] fourth_order_double_sin_cos_K1_q0;
    wire   [7:0] fourth_order_double_sin_cos_K2_address0;
    reg    fourth_order_double_sin_cos_K2_ce0;
    wire   [43:0] fourth_order_double_sin_cos_K2_q0;
    wire   [7:0] fourth_order_double_sin_cos_K3_address0;
    reg    fourth_order_double_sin_cos_K3_ce0;
    wire   [32:0] fourth_order_double_sin_cos_K3_q0;
    wire   [7:0] fourth_order_double_sin_cos_K4_address0;
    reg    fourth_order_double_sin_cos_K4_ce0;
    wire   [24:0] fourth_order_double_sin_cos_K4_q0;
    reg   [0:0] do_cos_read_reg_1592;
    wire    ap_block_pp0_stage0_11001;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter1_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter2_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter3_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter4_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter5_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter6_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter7_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter8_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter9_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter10_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter11_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter12_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter13_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter14_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter15_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter16_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter17_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter18_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter19_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter20_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter21_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter22_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter23_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter24_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter25_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter26_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter27_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter28_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter29_reg;
    reg   [0:0] do_cos_read_reg_1592_pp0_iter30_reg;
    reg   [0:0] din_sign_reg_1600;
    reg   [0:0] din_sign_reg_1600_pp0_iter1_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter2_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter3_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter4_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter5_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter6_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter7_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter8_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter9_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter10_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter11_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter12_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter13_reg;
    reg   [0:0] din_sign_reg_1600_pp0_iter14_reg;
    wire   [10:0] din_exp_fu_396_p4;
    reg   [10:0] din_exp_reg_1606;
    reg   [10:0] din_exp_reg_1606_pp0_iter1_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter2_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter3_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter4_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter5_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter6_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter7_reg;
    reg   [10:0] din_exp_reg_1606_pp0_iter8_reg;
    wire   [51:0] din_sig_fu_406_p1;
    reg   [51:0] din_sig_reg_1613;
    reg   [51:0] din_sig_reg_1613_pp0_iter1_reg;
    reg   [51:0] din_sig_reg_1613_pp0_iter2_reg;
    wire   [0:0] closepath_fu_410_p2;
    reg   [0:0] closepath_reg_1619;
    reg   [0:0] closepath_reg_1619_pp0_iter1_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter2_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter3_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter4_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter5_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter6_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter7_reg;
    reg   [0:0] closepath_reg_1619_pp0_iter8_reg;
    wire   [6:0] trunc_ln398_fu_445_p1;
    reg   [6:0] trunc_ln398_reg_1631;
    reg   [6:0] trunc_ln398_reg_1631_pp0_iter1_reg;
    reg   [255:0] table_256_reg_1636;
    reg  signed [169:0] Med_reg_1641;
    wire   [0:0] icmp_ln271_1_fu_479_p2;
    reg   [0:0] icmp_ln271_1_reg_1651;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter4_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter5_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter6_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter7_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter8_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter9_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter10_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter11_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter12_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter13_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter14_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter15_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter16_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter17_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter18_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter19_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter20_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter21_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter22_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter23_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter24_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter25_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter26_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter27_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter28_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter29_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter30_reg;
    reg   [0:0] icmp_ln271_1_reg_1651_pp0_iter31_reg;
    wire   [169:0] grp_fu_380_p2;
    reg   [169:0] h_reg_1657;
    reg   [123:0] Mx_bits_reg_1662;
    reg   [2:0] k_reg_1668;
    reg   [2:0] k_reg_1668_pp0_iter8_reg;
    wire   [123:0] Mx_bits_3_fu_527_p3;
    reg   [123:0] Mx_bits_3_reg_1673;
    wire   [6:0] Mx_zeros_fu_582_p1;
    reg   [6:0] Mx_zeros_reg_1678;
    wire   [2:0] k_1_fu_598_p3;
    reg   [2:0] k_1_reg_1684;
    reg   [2:0] k_1_reg_1684_pp0_iter10_reg;
    reg   [2:0] k_1_reg_1684_pp0_iter11_reg;
    reg   [2:0] k_1_reg_1684_pp0_iter12_reg;
    reg   [2:0] k_1_reg_1684_pp0_iter13_reg;
    reg   [62:0] Mx_reg_1690;
    reg   [62:0] Mx_reg_1690_pp0_iter10_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter11_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter12_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter13_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter14_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter15_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter16_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter17_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter18_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter19_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter20_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter21_reg;
    reg   [62:0] Mx_reg_1690_pp0_iter22_reg;
    wire   [10:0] Ex_1_fu_625_p2;
    reg   [10:0] Ex_1_reg_1697;
    reg   [10:0] Ex_1_reg_1697_pp0_iter10_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter11_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter12_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter13_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter14_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter15_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter16_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter17_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter18_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter19_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter20_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter21_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter22_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter23_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter24_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter25_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter26_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter27_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter28_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter29_reg;
    reg   [10:0] Ex_1_reg_1697_pp0_iter30_reg;
    reg   [0:0] tmp_3_reg_1703;
    wire   [10:0] sub_ln506_fu_639_p2;
    reg   [10:0] sub_ln506_reg_1709;
    wire   [0:0] icmp_ln271_fu_645_p2;
    reg   [0:0] icmp_ln271_reg_1714;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter10_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter11_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter12_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter13_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter14_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter15_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter16_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter17_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter18_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter19_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter20_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter21_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter22_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter23_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter24_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter25_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter26_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter27_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter28_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter29_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter30_reg;
    reg   [0:0] icmp_ln271_reg_1714_pp0_iter31_reg;
    wire   [0:0] icmp_ln282_fu_650_p2;
    reg   [0:0] icmp_ln282_reg_1720;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter10_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter11_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter12_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter13_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter14_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter15_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter16_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter17_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter18_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter19_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter20_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter21_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter22_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter23_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter24_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter25_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter26_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter27_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter28_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter29_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter30_reg;
    reg   [0:0] icmp_ln282_reg_1720_pp0_iter31_reg;
    reg   [6:0] tmp_8_reg_1728;
    reg   [6:0] tmp_8_reg_1728_pp0_iter11_reg;
    reg   [6:0] tmp_8_reg_1728_pp0_iter12_reg;
    reg   [6:0] tmp_8_reg_1728_pp0_iter13_reg;
    wire   [55:0] B_fu_691_p1;
    reg   [55:0] B_reg_1733;
    reg   [55:0] B_reg_1733_pp0_iter11_reg;
    reg   [55:0] B_reg_1733_pp0_iter12_reg;
    reg   [55:0] B_reg_1733_pp0_iter13_reg;
    reg   [55:0] B_reg_1733_pp0_iter14_reg;
    reg   [55:0] B_reg_1733_pp0_iter15_reg;
    reg   [48:0] B_trunc_reg_1738;
    wire   [97:0] zext_ln25_fu_705_p1;
    reg   [97:0] zext_ln25_reg_1743;
    reg   [97:0] zext_ln25_reg_1743_pp0_iter12_reg;
    reg   [97:0] zext_ln25_reg_1743_pp0_iter13_reg;
    reg   [97:0] zext_ln25_reg_1743_pp0_iter14_reg;
    reg   [97:0] zext_ln25_reg_1743_pp0_iter15_reg;
    wire   [0:0] cos_basis_fu_755_p3;
    reg   [0:0] cos_basis_reg_1750;
    reg   [0:0] cos_basis_reg_1750_pp0_iter15_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter16_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter17_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter18_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter19_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter20_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter21_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter22_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter23_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter24_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter25_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter26_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter27_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter28_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter29_reg;
    reg   [0:0] cos_basis_reg_1750_pp0_iter30_reg;
    wire   [63:0] zext_ln32_fu_776_p1;
    reg   [63:0] zext_ln32_reg_1756;
    reg   [63:0] zext_ln32_reg_1756_pp0_iter15_reg;
    reg   [63:0] zext_ln32_reg_1756_pp0_iter16_reg;
    reg   [63:0] zext_ln32_reg_1756_pp0_iter17_reg;
    reg   [63:0] zext_ln32_reg_1756_pp0_iter18_reg;
    wire   [0:0] results_sign_3_fu_945_p2;
    reg   [0:0] results_sign_3_reg_1773;
    reg   [48:0] B_squared_reg_1778;
    reg  signed [51:0] fourth_order_double_sin_cos_K1_load_reg_1784;
    reg  signed [43:0] fourth_order_double_sin_cos_K2_load_reg_1789;
    wire   [0:0] and_ln271_fu_961_p2;
    reg   [0:0] and_ln271_reg_1794;
    reg   [0:0] and_ln271_reg_1794_pp0_iter16_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter17_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter18_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter19_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter20_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter21_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter22_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter23_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter24_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter25_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter26_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter27_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter28_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter29_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter30_reg;
    reg   [0:0] and_ln271_reg_1794_pp0_iter31_reg;
    wire   [0:0] results_sign_4_fu_975_p3;
    reg   [0:0] results_sign_4_reg_1800;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter16_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter17_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter18_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter19_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter20_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter21_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter22_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter23_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter24_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter25_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter26_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter27_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter28_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter29_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter30_reg;
    reg   [0:0] results_sign_4_reg_1800_pp0_iter31_reg;
    wire   [97:0] zext_ln25_1_fu_982_p1;
    reg   [58:0] t1_reg_1847;
    reg   [55:0] trunc_ln_reg_1852;
    reg   [47:0] trunc_ln1_reg_1857;
    reg   [41:0] tmp_10_reg_1862;
    reg   [32:0] fourth_order_double_sin_cos_K3_load_reg_1867;
    reg   [34:0] tmp_11_reg_1872;
    reg   [24:0] fourth_order_double_sin_cos_K4_load_reg_1877;
    wire   [63:0] add_ln37_1_fu_1083_p2;
    reg   [63:0] add_ln37_1_reg_1902;
    reg   [63:0] add_ln37_1_reg_1902_pp0_iter22_reg;
    reg   [28:0] lshr_ln_reg_1907;
    reg   [36:0] tmp_12_reg_1912;
    wire   [62:0] Mx_1_fu_1109_p3;
    reg   [62:0] Mx_1_reg_1917;
    wire   [63:0] add_ln37_3_fu_1126_p2;
    reg  signed [63:0] add_ln37_3_reg_1922;
    reg   [62:0] result_reg_1937;
    reg   [15:0] tmp_i_reg_1943;
    reg   [15:0] tmp_3_i_reg_1948;
    reg   [15:0] tmp_3_i_reg_1948_pp0_iter29_reg;
    reg   [15:0] tmp_6_i_reg_1953;
    reg   [15:0] tmp_6_i_reg_1953_pp0_iter29_reg;
    reg   [14:0] tmp_9_i_reg_1958;
    reg   [14:0] tmp_9_i_reg_1958_pp0_iter29_reg;
    reg   [14:0] tmp_9_i_reg_1958_pp0_iter30_reg;
    reg   [31:0] c_fu_1207_p3;
    reg   [31:0] c_reg_1963;
    reg   [31:0] c_reg_1963_pp0_iter30_reg;
    wire   [62:0] in_shift_1_fu_1219_p2;
    reg   [62:0] in_shift_1_reg_1969;
    reg   [62:0] in_shift_1_reg_1969_pp0_iter30_reg;
    wire   [0:0] icmp_ln433_fu_1224_p2;
    reg   [0:0] icmp_ln433_reg_1975;
    reg   [0:0] icmp_ln433_reg_1975_pp0_iter30_reg;
    reg   [31:0] c_2_fu_1271_p3;
    reg   [31:0] c_2_reg_1980;
    wire   [0:0] icmp_ln424_fu_1279_p2;
    reg   [0:0] icmp_ln424_reg_1985;
    wire   [31:0] shift_1_fu_1284_p2;
    reg   [31:0] shift_1_reg_1993;
    wire   [62:0] in_shift_2_fu_1294_p2;
    reg   [62:0] in_shift_2_reg_1998;
    reg   [62:0] in_shift_2_reg_1998_pp0_iter31_reg;
    wire   [0:0] icmp_ln424_1_fu_1299_p2;
    reg   [0:0] icmp_ln424_1_reg_2004;
    wire   [31:0] shift_2_fu_1305_p2;
    reg   [31:0] shift_2_reg_2010;
    wire   [0:0] icmp_ln424_2_fu_1311_p2;
    reg   [0:0] icmp_ln424_2_reg_2016;
    reg   [31:0] c_3_fu_1344_p3;
    reg   [31:0] c_3_reg_2021;
    wire   [62:0] in_shift_3_fu_1355_p2;
    reg   [62:0] in_shift_3_reg_2026;
    wire   [0:0] and_ln424_2_fu_1379_p2;
    reg   [0:0] and_ln424_2_reg_2031;
    wire   [0:0] or_ln424_fu_1391_p2;
    reg   [0:0] or_ln424_reg_2036;
    wire   [0:0] or_ln433_fu_1434_p2;
    reg   [0:0] or_ln433_reg_2041;
    wire   [51:0] select_ln424_4_fu_1458_p3;
    reg   [51:0] select_ln424_4_reg_2046;
    wire   [10:0] results_exp_1_fu_1496_p3;
    reg   [10:0] results_exp_1_reg_2051;
    wire   [63:0] zext_ln397_fu_440_p1;
    wire    ap_block_pp0_stage0;
    wire   [34:0] grp_fu_348_p0;
    wire   [24:0] grp_fu_348_p1;
    wire   [41:0] grp_fu_352_p0;
    wire   [32:0] grp_fu_352_p1;
    wire   [48:0] grp_fu_356_p0;
    wire   [48:0] grp_fu_360_p0;
    wire   [48:0] grp_fu_360_p1;
    wire   [48:0] grp_fu_364_p0;
    wire   [48:0] grp_fu_364_p1;
    wire   [48:0] grp_fu_368_p0;
    wire   [48:0] grp_fu_368_p1;
    wire   [55:0] grp_fu_372_p0;
    wire   [62:0] grp_fu_376_p1;
    wire   [52:0] grp_fu_380_p1;
    wire   [63:0] data_fu_384_p1;
    wire   [10:0] add_ln396_fu_416_p2;
    wire   [10:0] addr_fu_422_p3;
    wire   [3:0] tmp_s_fu_430_p4;
    wire   [255:0] zext_ln398_fu_449_p1;
    wire   [255:0] shl_ln398_fu_452_p2;
    wire   [52:0] X_fu_467_p3;
    wire   [0:0] tmp_fu_504_p3;
    wire   [0:0] xor_ln451_fu_511_p2;
    wire   [0:0] and_ln451_fu_516_p2;
    wire   [123:0] Mx_bits_1_fu_522_p2;
    wire   [60:0] tmp_1_fu_534_p4;
    wire   [61:0] t_fu_544_p3;
    reg   [61:0] tmp_4_fu_552_p4;
    wire   [62:0] tmp_5_fu_562_p3;
    wire  signed [63:0] sext_ln75_fu_570_p1;
    reg   [63:0] tmp_6_fu_574_p3;
    wire   [10:0] Ex_fu_586_p2;
    wire   [123:0] zext_ln504_fu_607_p1;
    wire   [123:0] shl_ln504_fu_610_p2;
    wire   [10:0] select_ln453_fu_591_p3;
    wire   [10:0] zext_ln505_fu_604_p1;
    wire   [10:0] select_ln506_fu_655_p3;
    wire   [62:0] zext_ln506_fu_660_p1;
    wire   [62:0] lshr_ln506_fu_664_p2;
    wire   [62:0] shl_ln506_fu_669_p2;
    wire   [62:0] x_1_fu_674_p3;
    wire   [0:0] tmp_7_fu_710_p17;
    wire   [0:0] tmp_7_fu_710_p19;
    wire   [0:0] xor_ln242_fu_749_p2;
    wire   [0:0] sin_basis_fu_762_p3;
    wire   [7:0] A_fu_769_p3;
    wire   [0:0] tmp_9_fu_788_p33;
    wire   [3:0] index_fu_782_p3;
    wire   [0:0] tmp_2_fu_860_p33;
    wire   [0:0] tmp_9_fu_788_p35;
    wire   [0:0] tmp_2_fu_860_p35;
    wire   [0:0] results_sign_fu_932_p3;
    wire   [0:0] xor_ln282_fu_940_p2;
    wire   [97:0] grp_fu_360_p2;
    wire   [0:0] xor_ln278_fu_965_p2;
    wire   [0:0] results_sign_2_fu_970_p2;
    wire   [107:0] grp_fu_372_p2;
    wire   [92:0] grp_fu_356_p2;
    wire   [97:0] grp_fu_364_p2;
    wire   [97:0] grp_fu_368_p2;
    wire   [62:0] t1_1_fu_1044_p3;
    wire  signed [63:0] sext_ln37_fu_1067_p1;
    wire  signed [63:0] sext_ln37_1_fu_1071_p1;
    wire   [63:0] add_ln37_fu_1074_p2;
    wire  signed [63:0] sext_ln37_2_fu_1080_p1;
    wire   [59:0] grp_fu_348_p2;
    wire   [74:0] grp_fu_352_p2;
    wire   [63:0] zext_ln37_2_fu_1115_p1;
    wire   [63:0] add_ln37_2_fu_1118_p2;
    wire   [63:0] zext_ln37_fu_1123_p1;
    wire   [125:0] grp_fu_376_p2;
    wire   [31:0] out_bits_fu_1190_p3;
    reg   [31:0] tmp_2_i_fu_1197_p4;
    wire   [62:0] zext_ln423_fu_1215_p1;
    wire   [31:0] out_bits_4_fu_1229_p3;
    reg   [31:0] tmp_5_i_fu_1243_p4;
    wire   [31:0] out_bits_5_fu_1236_p3;
    reg   [31:0] tmp_8_i_fu_1261_p4;
    reg   [31:0] c_1_fu_1253_p3;
    wire   [62:0] zext_ln423_1_fu_1290_p1;
    wire   [10:0] Ex_2_fu_1317_p3;
    wire   [31:0] out_bits_6_fu_1327_p3;
    reg   [31:0] tmp_i_63_fu_1334_p4;
    wire   [62:0] zext_ln423_2_fu_1352_p1;
    wire   [0:0] and_ln424_fu_1365_p2;
    wire   [0:0] xor_ln424_fu_1374_p2;
    wire   [31:0] add_ln422_fu_1360_p2;
    wire   [0:0] and_ln424_1_fu_1369_p2;
    wire   [31:0] select_ln424_fu_1384_p3;
    wire   [31:0] select_ln424_1_fu_1397_p3;
    wire  signed [11:0] sext_ln252_fu_1323_p1;
    wire   [11:0] add_ln432_fu_1410_p2;
    wire  signed [31:0] sext_ln432_fu_1416_p1;
    wire   [31:0] select_ln424_2_fu_1402_p3;
    wire   [31:0] newexp_fu_1420_p2;
    wire   [0:0] tmp_13_fu_1426_p3;
    wire   [51:0] tmp_16_fu_1439_p4;
    wire   [51:0] tmp_17_fu_1449_p4;
    wire   [0:0] or_ln282_fu_1483_p2;
    wire   [10:0] select_ln282_fu_1476_p3;
    wire   [10:0] empty_fu_1465_p1;
    wire   [10:0] select_ln259_fu_1469_p3;
    wire   [10:0] results_exp_fu_1488_p3;
    wire   [62:0] zext_ln423_3_fu_1503_p1;
    wire   [62:0] shl_ln423_fu_1506_p2;
    wire   [51:0] tmp_14_fu_1511_p4;
    wire   [51:0] tmp_15_fu_1520_p4;
    wire   [51:0] select_ln424_3_fu_1530_p3;
    wire   [51:0] select_ln424_5_fu_1537_p3;
    wire   [0:0] and_ln271_1_fu_1550_p2;
    wire   [0:0] xor_ln271_fu_1554_p2;
    wire   [0:0] or_ln271_fu_1568_p2;
    wire   [51:0] select_ln271_fu_1560_p3;
    wire   [51:0] significand_fu_1543_p3;
    wire   [51:0] results_sig_1_fu_1572_p3;
    wire   [63:0] t_2_fu_1580_p4;
    reg    grp_fu_348_ce;
    reg    grp_fu_352_ce;
    reg    grp_fu_356_ce;
    reg    grp_fu_360_ce;
    reg    grp_fu_364_ce;
    reg    grp_fu_368_ce;
    reg    grp_fu_372_ce;
    reg    grp_fu_376_ce;
    reg    grp_fu_380_ce;
    reg   [0:0] ap_NS_fsm;
    reg    ap_idle_pp0_0to31;
    reg    ap_reset_idle_pp0;
    wire    ap_enable_pp0;
    wire   [59:0] grp_fu_348_p00;
    wire   [59:0] grp_fu_348_p10;
    wire   [74:0] grp_fu_352_p00;
    wire   [74:0] grp_fu_352_p10;
    wire   [92:0] grp_fu_356_p00;
    wire   [107:0] grp_fu_372_p00;
    wire   [125:0] grp_fu_376_p10;
    wire   [169:0] grp_fu_380_p10;
    wire   [2:0] tmp_7_fu_710_p1;
    wire   [2:0] tmp_7_fu_710_p3;
    wire   [2:0] tmp_7_fu_710_p5;
    wire   [2:0] tmp_7_fu_710_p7;
    wire  signed [2:0] tmp_7_fu_710_p9;
    wire  signed [2:0] tmp_7_fu_710_p11;
    wire  signed [2:0] tmp_7_fu_710_p13;
    wire  signed [2:0] tmp_7_fu_710_p15;
    wire   [3:0] tmp_9_fu_788_p1;
    wire   [3:0] tmp_9_fu_788_p3;
    wire   [3:0] tmp_9_fu_788_p5;
    wire   [3:0] tmp_9_fu_788_p7;
    wire   [3:0] tmp_9_fu_788_p9;
    wire   [3:0] tmp_9_fu_788_p11;
    wire   [3:0] tmp_9_fu_788_p13;
    wire   [3:0] tmp_9_fu_788_p15;
    wire  signed [3:0] tmp_9_fu_788_p17;
    wire  signed [3:0] tmp_9_fu_788_p19;
    wire  signed [3:0] tmp_9_fu_788_p21;
    wire  signed [3:0] tmp_9_fu_788_p23;
    wire  signed [3:0] tmp_9_fu_788_p25;
    wire  signed [3:0] tmp_9_fu_788_p27;
    wire  signed [3:0] tmp_9_fu_788_p29;
    wire  signed [3:0] tmp_9_fu_788_p31;
    wire   [3:0] tmp_2_fu_860_p1;
    wire   [3:0] tmp_2_fu_860_p3;
    wire   [3:0] tmp_2_fu_860_p5;
    wire   [3:0] tmp_2_fu_860_p7;
    wire   [3:0] tmp_2_fu_860_p9;
    wire   [3:0] tmp_2_fu_860_p11;
    wire   [3:0] tmp_2_fu_860_p13;
    wire   [3:0] tmp_2_fu_860_p15;
    wire  signed [3:0] tmp_2_fu_860_p17;
    wire  signed [3:0] tmp_2_fu_860_p19;
    wire  signed [3:0] tmp_2_fu_860_p21;
    wire  signed [3:0] tmp_2_fu_860_p23;
    wire  signed [3:0] tmp_2_fu_860_p25;
    wire  signed [3:0] tmp_2_fu_860_p27;
    wire  signed [3:0] tmp_2_fu_860_p29;
    wire  signed [3:0] tmp_2_fu_860_p31;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 1'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter10 = 1'b0;
        #0 ap_enable_reg_pp0_iter11 = 1'b0;
        #0 ap_enable_reg_pp0_iter12 = 1'b0;
        #0 ap_enable_reg_pp0_iter13 = 1'b0;
        #0 ap_enable_reg_pp0_iter14 = 1'b0;
        #0 ap_enable_reg_pp0_iter15 = 1'b0;
        #0 ap_enable_reg_pp0_iter16 = 1'b0;
        #0 ap_enable_reg_pp0_iter17 = 1'b0;
        #0 ap_enable_reg_pp0_iter18 = 1'b0;
        #0 ap_enable_reg_pp0_iter19 = 1'b0;
        #0 ap_enable_reg_pp0_iter20 = 1'b0;
        #0 ap_enable_reg_pp0_iter21 = 1'b0;
        #0 ap_enable_reg_pp0_iter22 = 1'b0;
        #0 ap_enable_reg_pp0_iter23 = 1'b0;
        #0 ap_enable_reg_pp0_iter24 = 1'b0;
        #0 ap_enable_reg_pp0_iter25 = 1'b0;
        #0 ap_enable_reg_pp0_iter26 = 1'b0;
        #0 ap_enable_reg_pp0_iter27 = 1'b0;
        #0 ap_enable_reg_pp0_iter28 = 1'b0;
        #0 ap_enable_reg_pp0_iter29 = 1'b0;
        #0 ap_enable_reg_pp0_iter30 = 1'b0;
        #0 ap_enable_reg_pp0_iter31 = 1'b0;
        #0 ap_enable_reg_pp0_iter32 = 1'b0;
    end

    main_sin_or_cos_double_s_ref_4oPi_table_256_ROM_AUTO_1R #(
        .DataWidth(256),
        .AddressRange(10),
        .AddressWidth(4)
    ) ref_4oPi_table_256_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(ref_4oPi_table_256_address0),
        .ce0(ref_4oPi_table_256_ce0),
        .q0(ref_4oPi_table_256_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K0_ROM_1P_LUTRAM_1R #(
        .DataWidth(59),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K0_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K0_address0),
        .ce0(fourth_order_double_sin_cos_K0_ce0),
        .q0(fourth_order_double_sin_cos_K0_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K1_ROM_1P_LUTRAM_1R #(
        .DataWidth(52),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K1_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K1_address0),
        .ce0(fourth_order_double_sin_cos_K1_ce0),
        .q0(fourth_order_double_sin_cos_K1_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K2_ROM_1P_LUTRAM_1R #(
        .DataWidth(44),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K2_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K2_address0),
        .ce0(fourth_order_double_sin_cos_K2_ce0),
        .q0(fourth_order_double_sin_cos_K2_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K3_ROM_1P_LUTRAM_1R #(
        .DataWidth(33),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K3_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K3_address0),
        .ce0(fourth_order_double_sin_cos_K3_ce0),
        .q0(fourth_order_double_sin_cos_K3_q0)
    );

    main_sin_or_cos_double_s_fourth_order_double_sin_cos_K4_ROM_1P_LUTRAM_1R #(
        .DataWidth(25),
        .AddressRange(256),
        .AddressWidth(8)
    ) fourth_order_double_sin_cos_K4_U (
        .clk(ap_clk),
        .reset(ap_rst),
        .address0(fourth_order_double_sin_cos_K4_address0),
        .ce0(fourth_order_double_sin_cos_K4_ce0),
        .q0(fourth_order_double_sin_cos_K4_q0)
    );

    main_mul_35ns_25ns_60_2_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(35),
        .din1_WIDTH(25),
        .dout_WIDTH(60)
    ) mul_35ns_25ns_60_2_1_U345 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_348_p0),
        .din1(grp_fu_348_p1),
        .ce(grp_fu_348_ce),
        .dout(grp_fu_348_p2)
    );

    main_mul_42ns_33ns_75_2_1 #(
        .ID(1),
        .NUM_STAGE(2),
        .din0_WIDTH(42),
        .din1_WIDTH(33),
        .dout_WIDTH(75)
    ) mul_42ns_33ns_75_2_1_U346 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_352_p0),
        .din1(grp_fu_352_p1),
        .ce(grp_fu_352_ce),
        .dout(grp_fu_352_p2)
    );

    main_mul_49ns_44s_93_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(44),
        .dout_WIDTH(93)
    ) mul_49ns_44s_93_5_1_U347 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_356_p0),
        .din1(fourth_order_double_sin_cos_K2_load_reg_1789),
        .ce(grp_fu_356_ce),
        .dout(grp_fu_356_p2)
    );

    main_mul_49ns_49ns_98_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(49),
        .dout_WIDTH(98)
    ) mul_49ns_49ns_98_5_1_U348 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_360_p0),
        .din1(grp_fu_360_p1),
        .ce(grp_fu_360_ce),
        .dout(grp_fu_360_p2)
    );

    main_mul_49ns_49ns_98_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(49),
        .dout_WIDTH(98)
    ) mul_49ns_49ns_98_5_1_U349 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_364_p0),
        .din1(grp_fu_364_p1),
        .ce(grp_fu_364_ce),
        .dout(grp_fu_364_p2)
    );

    main_mul_49ns_49ns_98_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(49),
        .din1_WIDTH(49),
        .dout_WIDTH(98)
    ) mul_49ns_49ns_98_5_1_U350 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_368_p0),
        .din1(grp_fu_368_p1),
        .ce(grp_fu_368_ce),
        .dout(grp_fu_368_p2)
    );

    main_mul_56ns_52s_108_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(56),
        .din1_WIDTH(52),
        .dout_WIDTH(108)
    ) mul_56ns_52s_108_5_1_U351 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_372_p0),
        .din1(fourth_order_double_sin_cos_K1_load_reg_1784),
        .ce(grp_fu_372_ce),
        .dout(grp_fu_372_p2)
    );

    main_mul_64s_63ns_126_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(64),
        .din1_WIDTH(63),
        .dout_WIDTH(126)
    ) mul_64s_63ns_126_5_1_U352 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(add_ln37_3_reg_1922),
        .din1(grp_fu_376_p1),
        .ce(grp_fu_376_ce),
        .dout(grp_fu_376_p2)
    );

    main_mul_170s_53ns_170_5_1 #(
        .ID(1),
        .NUM_STAGE(5),
        .din0_WIDTH(170),
        .din1_WIDTH(53),
        .dout_WIDTH(170)
    ) mul_170s_53ns_170_5_1_U353 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(Med_reg_1641),
        .din1(grp_fu_380_p1),
        .ce(grp_fu_380_ce),
        .dout(grp_fu_380_p2)
    );

    main_sparsemux_17_3_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(3'h0),
        .din0_WIDTH(1),
        .CASE1(3'h1),
        .din1_WIDTH(1),
        .CASE2(3'h2),
        .din2_WIDTH(1),
        .CASE3(3'h3),
        .din3_WIDTH(1),
        .CASE4(3'h4),
        .din4_WIDTH(1),
        .CASE5(3'h5),
        .din5_WIDTH(1),
        .CASE6(3'h6),
        .din6_WIDTH(1),
        .CASE7(3'h7),
        .din7_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(3),
        .dout_WIDTH(1)
    ) sparsemux_17_3_1_1_1_U354 (
        .din0(1'd0),
        .din1(1'd1),
        .din2(1'd1),
        .din3(1'd0),
        .din4(1'd0),
        .din5(1'd1),
        .din6(1'd1),
        .din7(1'd0),
        .def (tmp_7_fu_710_p17),
        .sel (k_1_reg_1684_pp0_iter13_reg),
        .dout(tmp_7_fu_710_p19)
    );

    main_sparsemux_33_4_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(4'h0),
        .din0_WIDTH(1),
        .CASE1(4'h1),
        .din1_WIDTH(1),
        .CASE2(4'h2),
        .din2_WIDTH(1),
        .CASE3(4'h3),
        .din3_WIDTH(1),
        .CASE4(4'h4),
        .din4_WIDTH(1),
        .CASE5(4'h5),
        .din5_WIDTH(1),
        .CASE6(4'h6),
        .din6_WIDTH(1),
        .CASE7(4'h7),
        .din7_WIDTH(1),
        .CASE8(4'h8),
        .din8_WIDTH(1),
        .CASE9(4'h9),
        .din9_WIDTH(1),
        .CASE10(4'hA),
        .din10_WIDTH(1),
        .CASE11(4'hB),
        .din11_WIDTH(1),
        .CASE12(4'hC),
        .din12_WIDTH(1),
        .CASE13(4'hD),
        .din13_WIDTH(1),
        .CASE14(4'hE),
        .din14_WIDTH(1),
        .CASE15(4'hF),
        .din15_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(4),
        .dout_WIDTH(1)
    ) sparsemux_33_4_1_1_1_U355 (
        .din0 (1'd0),
        .din1 (1'd0),
        .din2 (1'd0),
        .din3 (1'd1),
        .din4 (1'd1),
        .din5 (1'd1),
        .din6 (1'd1),
        .din7 (1'd0),
        .din8 (1'd0),
        .din9 (1'd1),
        .din10(1'd1),
        .din11(1'd1),
        .din12(1'd1),
        .din13(1'd0),
        .din14(1'd0),
        .din15(1'd0),
        .def  (tmp_9_fu_788_p33),
        .sel  (index_fu_782_p3),
        .dout (tmp_9_fu_788_p35)
    );

    main_sparsemux_33_4_1_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .CASE0(4'h0),
        .din0_WIDTH(1),
        .CASE1(4'h1),
        .din1_WIDTH(1),
        .CASE2(4'h2),
        .din2_WIDTH(1),
        .CASE3(4'h3),
        .din3_WIDTH(1),
        .CASE4(4'h4),
        .din4_WIDTH(1),
        .CASE5(4'h5),
        .din5_WIDTH(1),
        .CASE6(4'h6),
        .din6_WIDTH(1),
        .CASE7(4'h7),
        .din7_WIDTH(1),
        .CASE8(4'h8),
        .din8_WIDTH(1),
        .CASE9(4'h9),
        .din9_WIDTH(1),
        .CASE10(4'hA),
        .din10_WIDTH(1),
        .CASE11(4'hB),
        .din11_WIDTH(1),
        .CASE12(4'hC),
        .din12_WIDTH(1),
        .CASE13(4'hD),
        .din13_WIDTH(1),
        .CASE14(4'hE),
        .din14_WIDTH(1),
        .CASE15(4'hF),
        .din15_WIDTH(1),
        .def_WIDTH(1),
        .sel_WIDTH(4),
        .dout_WIDTH(1)
    ) sparsemux_33_4_1_1_1_U356 (
        .din0 (1'd0),
        .din1 (1'd0),
        .din2 (1'd1),
        .din3 (1'd0),
        .din4 (1'd1),
        .din5 (1'd1),
        .din6 (1'd0),
        .din7 (1'd1),
        .din8 (1'd1),
        .din9 (1'd0),
        .din10(1'd1),
        .din11(1'd1),
        .din12(1'd0),
        .din13(1'd1),
        .din14(1'd0),
        .din15(1'd0),
        .def  (tmp_2_fu_860_p33),
        .sel  (index_fu_782_p3),
        .dout (tmp_2_fu_860_p35)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_enable_reg_pp0_iter1 <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter10 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter11 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter12 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter13 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter14 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter15 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter16 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter17 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter18 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter19 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter20 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter21 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter23 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter23 <= ap_enable_reg_pp0_iter22;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter24 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter24 <= ap_enable_reg_pp0_iter23;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter25 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter25 <= ap_enable_reg_pp0_iter24;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter26 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter26 <= ap_enable_reg_pp0_iter25;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter27 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter27 <= ap_enable_reg_pp0_iter26;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter28 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter28 <= ap_enable_reg_pp0_iter27;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter29 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter29 <= ap_enable_reg_pp0_iter28;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter30 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter30 <= ap_enable_reg_pp0_iter29;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter31 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter31 <= ap_enable_reg_pp0_iter30;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter32 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter32 <= ap_enable_reg_pp0_iter31;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            B_reg_1733 <= B_fu_691_p1;
            B_reg_1733_pp0_iter11_reg <= B_reg_1733;
            B_reg_1733_pp0_iter12_reg <= B_reg_1733_pp0_iter11_reg;
            B_reg_1733_pp0_iter13_reg <= B_reg_1733_pp0_iter12_reg;
            B_reg_1733_pp0_iter14_reg <= B_reg_1733_pp0_iter13_reg;
            B_reg_1733_pp0_iter15_reg <= B_reg_1733_pp0_iter14_reg;
            B_squared_reg_1778 <= {{grp_fu_360_p2[97:49]}};
            B_trunc_reg_1738 <= {{x_1_fu_674_p3[55:7]}};
            Ex_1_reg_1697 <= Ex_1_fu_625_p2;
            Ex_1_reg_1697_pp0_iter10_reg <= Ex_1_reg_1697;
            Ex_1_reg_1697_pp0_iter11_reg <= Ex_1_reg_1697_pp0_iter10_reg;
            Ex_1_reg_1697_pp0_iter12_reg <= Ex_1_reg_1697_pp0_iter11_reg;
            Ex_1_reg_1697_pp0_iter13_reg <= Ex_1_reg_1697_pp0_iter12_reg;
            Ex_1_reg_1697_pp0_iter14_reg <= Ex_1_reg_1697_pp0_iter13_reg;
            Ex_1_reg_1697_pp0_iter15_reg <= Ex_1_reg_1697_pp0_iter14_reg;
            Ex_1_reg_1697_pp0_iter16_reg <= Ex_1_reg_1697_pp0_iter15_reg;
            Ex_1_reg_1697_pp0_iter17_reg <= Ex_1_reg_1697_pp0_iter16_reg;
            Ex_1_reg_1697_pp0_iter18_reg <= Ex_1_reg_1697_pp0_iter17_reg;
            Ex_1_reg_1697_pp0_iter19_reg <= Ex_1_reg_1697_pp0_iter18_reg;
            Ex_1_reg_1697_pp0_iter20_reg <= Ex_1_reg_1697_pp0_iter19_reg;
            Ex_1_reg_1697_pp0_iter21_reg <= Ex_1_reg_1697_pp0_iter20_reg;
            Ex_1_reg_1697_pp0_iter22_reg <= Ex_1_reg_1697_pp0_iter21_reg;
            Ex_1_reg_1697_pp0_iter23_reg <= Ex_1_reg_1697_pp0_iter22_reg;
            Ex_1_reg_1697_pp0_iter24_reg <= Ex_1_reg_1697_pp0_iter23_reg;
            Ex_1_reg_1697_pp0_iter25_reg <= Ex_1_reg_1697_pp0_iter24_reg;
            Ex_1_reg_1697_pp0_iter26_reg <= Ex_1_reg_1697_pp0_iter25_reg;
            Ex_1_reg_1697_pp0_iter27_reg <= Ex_1_reg_1697_pp0_iter26_reg;
            Ex_1_reg_1697_pp0_iter28_reg <= Ex_1_reg_1697_pp0_iter27_reg;
            Ex_1_reg_1697_pp0_iter29_reg <= Ex_1_reg_1697_pp0_iter28_reg;
            Ex_1_reg_1697_pp0_iter30_reg <= Ex_1_reg_1697_pp0_iter29_reg;
            Med_reg_1641 <= {{shl_ln398_fu_452_p2[255:86]}};
            Mx_1_reg_1917 <= Mx_1_fu_1109_p3;
            Mx_bits_3_reg_1673 <= Mx_bits_3_fu_527_p3;
            Mx_bits_reg_1662 <= {{grp_fu_380_p2[166:43]}};
            Mx_reg_1690 <= {{shl_ln504_fu_610_p2[123:61]}};
            Mx_reg_1690_pp0_iter10_reg <= Mx_reg_1690;
            Mx_reg_1690_pp0_iter11_reg <= Mx_reg_1690_pp0_iter10_reg;
            Mx_reg_1690_pp0_iter12_reg <= Mx_reg_1690_pp0_iter11_reg;
            Mx_reg_1690_pp0_iter13_reg <= Mx_reg_1690_pp0_iter12_reg;
            Mx_reg_1690_pp0_iter14_reg <= Mx_reg_1690_pp0_iter13_reg;
            Mx_reg_1690_pp0_iter15_reg <= Mx_reg_1690_pp0_iter14_reg;
            Mx_reg_1690_pp0_iter16_reg <= Mx_reg_1690_pp0_iter15_reg;
            Mx_reg_1690_pp0_iter17_reg <= Mx_reg_1690_pp0_iter16_reg;
            Mx_reg_1690_pp0_iter18_reg <= Mx_reg_1690_pp0_iter17_reg;
            Mx_reg_1690_pp0_iter19_reg <= Mx_reg_1690_pp0_iter18_reg;
            Mx_reg_1690_pp0_iter20_reg <= Mx_reg_1690_pp0_iter19_reg;
            Mx_reg_1690_pp0_iter21_reg <= Mx_reg_1690_pp0_iter20_reg;
            Mx_reg_1690_pp0_iter22_reg <= Mx_reg_1690_pp0_iter21_reg;
            Mx_zeros_reg_1678 <= Mx_zeros_fu_582_p1;
            add_ln37_1_reg_1902 <= add_ln37_1_fu_1083_p2;
            add_ln37_1_reg_1902_pp0_iter22_reg <= add_ln37_1_reg_1902;
            add_ln37_3_reg_1922 <= add_ln37_3_fu_1126_p2;
            and_ln271_reg_1794 <= and_ln271_fu_961_p2;
            and_ln271_reg_1794_pp0_iter16_reg <= and_ln271_reg_1794;
            and_ln271_reg_1794_pp0_iter17_reg <= and_ln271_reg_1794_pp0_iter16_reg;
            and_ln271_reg_1794_pp0_iter18_reg <= and_ln271_reg_1794_pp0_iter17_reg;
            and_ln271_reg_1794_pp0_iter19_reg <= and_ln271_reg_1794_pp0_iter18_reg;
            and_ln271_reg_1794_pp0_iter20_reg <= and_ln271_reg_1794_pp0_iter19_reg;
            and_ln271_reg_1794_pp0_iter21_reg <= and_ln271_reg_1794_pp0_iter20_reg;
            and_ln271_reg_1794_pp0_iter22_reg <= and_ln271_reg_1794_pp0_iter21_reg;
            and_ln271_reg_1794_pp0_iter23_reg <= and_ln271_reg_1794_pp0_iter22_reg;
            and_ln271_reg_1794_pp0_iter24_reg <= and_ln271_reg_1794_pp0_iter23_reg;
            and_ln271_reg_1794_pp0_iter25_reg <= and_ln271_reg_1794_pp0_iter24_reg;
            and_ln271_reg_1794_pp0_iter26_reg <= and_ln271_reg_1794_pp0_iter25_reg;
            and_ln271_reg_1794_pp0_iter27_reg <= and_ln271_reg_1794_pp0_iter26_reg;
            and_ln271_reg_1794_pp0_iter28_reg <= and_ln271_reg_1794_pp0_iter27_reg;
            and_ln271_reg_1794_pp0_iter29_reg <= and_ln271_reg_1794_pp0_iter28_reg;
            and_ln271_reg_1794_pp0_iter30_reg <= and_ln271_reg_1794_pp0_iter29_reg;
            and_ln271_reg_1794_pp0_iter31_reg <= and_ln271_reg_1794_pp0_iter30_reg;
            and_ln424_2_reg_2031 <= and_ln424_2_fu_1379_p2;
            c_2_reg_1980 <= c_2_fu_1271_p3;
            c_3_reg_2021 <= c_3_fu_1344_p3;
            c_reg_1963 <= c_fu_1207_p3;
            c_reg_1963_pp0_iter30_reg <= c_reg_1963;
            closepath_reg_1619_pp0_iter2_reg <= closepath_reg_1619_pp0_iter1_reg;
            closepath_reg_1619_pp0_iter3_reg <= closepath_reg_1619_pp0_iter2_reg;
            closepath_reg_1619_pp0_iter4_reg <= closepath_reg_1619_pp0_iter3_reg;
            closepath_reg_1619_pp0_iter5_reg <= closepath_reg_1619_pp0_iter4_reg;
            closepath_reg_1619_pp0_iter6_reg <= closepath_reg_1619_pp0_iter5_reg;
            closepath_reg_1619_pp0_iter7_reg <= closepath_reg_1619_pp0_iter6_reg;
            closepath_reg_1619_pp0_iter8_reg <= closepath_reg_1619_pp0_iter7_reg;
            cos_basis_reg_1750 <= cos_basis_fu_755_p3;
            cos_basis_reg_1750_pp0_iter15_reg <= cos_basis_reg_1750;
            cos_basis_reg_1750_pp0_iter16_reg <= cos_basis_reg_1750_pp0_iter15_reg;
            cos_basis_reg_1750_pp0_iter17_reg <= cos_basis_reg_1750_pp0_iter16_reg;
            cos_basis_reg_1750_pp0_iter18_reg <= cos_basis_reg_1750_pp0_iter17_reg;
            cos_basis_reg_1750_pp0_iter19_reg <= cos_basis_reg_1750_pp0_iter18_reg;
            cos_basis_reg_1750_pp0_iter20_reg <= cos_basis_reg_1750_pp0_iter19_reg;
            cos_basis_reg_1750_pp0_iter21_reg <= cos_basis_reg_1750_pp0_iter20_reg;
            cos_basis_reg_1750_pp0_iter22_reg <= cos_basis_reg_1750_pp0_iter21_reg;
            cos_basis_reg_1750_pp0_iter23_reg <= cos_basis_reg_1750_pp0_iter22_reg;
            cos_basis_reg_1750_pp0_iter24_reg <= cos_basis_reg_1750_pp0_iter23_reg;
            cos_basis_reg_1750_pp0_iter25_reg <= cos_basis_reg_1750_pp0_iter24_reg;
            cos_basis_reg_1750_pp0_iter26_reg <= cos_basis_reg_1750_pp0_iter25_reg;
            cos_basis_reg_1750_pp0_iter27_reg <= cos_basis_reg_1750_pp0_iter26_reg;
            cos_basis_reg_1750_pp0_iter28_reg <= cos_basis_reg_1750_pp0_iter27_reg;
            cos_basis_reg_1750_pp0_iter29_reg <= cos_basis_reg_1750_pp0_iter28_reg;
            cos_basis_reg_1750_pp0_iter30_reg <= cos_basis_reg_1750_pp0_iter29_reg;
            din_exp_reg_1606_pp0_iter2_reg <= din_exp_reg_1606_pp0_iter1_reg;
            din_exp_reg_1606_pp0_iter3_reg <= din_exp_reg_1606_pp0_iter2_reg;
            din_exp_reg_1606_pp0_iter4_reg <= din_exp_reg_1606_pp0_iter3_reg;
            din_exp_reg_1606_pp0_iter5_reg <= din_exp_reg_1606_pp0_iter4_reg;
            din_exp_reg_1606_pp0_iter6_reg <= din_exp_reg_1606_pp0_iter5_reg;
            din_exp_reg_1606_pp0_iter7_reg <= din_exp_reg_1606_pp0_iter6_reg;
            din_exp_reg_1606_pp0_iter8_reg <= din_exp_reg_1606_pp0_iter7_reg;
            din_sig_reg_1613_pp0_iter2_reg <= din_sig_reg_1613_pp0_iter1_reg;
            din_sign_reg_1600_pp0_iter10_reg <= din_sign_reg_1600_pp0_iter9_reg;
            din_sign_reg_1600_pp0_iter11_reg <= din_sign_reg_1600_pp0_iter10_reg;
            din_sign_reg_1600_pp0_iter12_reg <= din_sign_reg_1600_pp0_iter11_reg;
            din_sign_reg_1600_pp0_iter13_reg <= din_sign_reg_1600_pp0_iter12_reg;
            din_sign_reg_1600_pp0_iter14_reg <= din_sign_reg_1600_pp0_iter13_reg;
            din_sign_reg_1600_pp0_iter2_reg <= din_sign_reg_1600_pp0_iter1_reg;
            din_sign_reg_1600_pp0_iter3_reg <= din_sign_reg_1600_pp0_iter2_reg;
            din_sign_reg_1600_pp0_iter4_reg <= din_sign_reg_1600_pp0_iter3_reg;
            din_sign_reg_1600_pp0_iter5_reg <= din_sign_reg_1600_pp0_iter4_reg;
            din_sign_reg_1600_pp0_iter6_reg <= din_sign_reg_1600_pp0_iter5_reg;
            din_sign_reg_1600_pp0_iter7_reg <= din_sign_reg_1600_pp0_iter6_reg;
            din_sign_reg_1600_pp0_iter8_reg <= din_sign_reg_1600_pp0_iter7_reg;
            din_sign_reg_1600_pp0_iter9_reg <= din_sign_reg_1600_pp0_iter8_reg;
            do_cos_read_reg_1592_pp0_iter10_reg <= do_cos_read_reg_1592_pp0_iter9_reg;
            do_cos_read_reg_1592_pp0_iter11_reg <= do_cos_read_reg_1592_pp0_iter10_reg;
            do_cos_read_reg_1592_pp0_iter12_reg <= do_cos_read_reg_1592_pp0_iter11_reg;
            do_cos_read_reg_1592_pp0_iter13_reg <= do_cos_read_reg_1592_pp0_iter12_reg;
            do_cos_read_reg_1592_pp0_iter14_reg <= do_cos_read_reg_1592_pp0_iter13_reg;
            do_cos_read_reg_1592_pp0_iter15_reg <= do_cos_read_reg_1592_pp0_iter14_reg;
            do_cos_read_reg_1592_pp0_iter16_reg <= do_cos_read_reg_1592_pp0_iter15_reg;
            do_cos_read_reg_1592_pp0_iter17_reg <= do_cos_read_reg_1592_pp0_iter16_reg;
            do_cos_read_reg_1592_pp0_iter18_reg <= do_cos_read_reg_1592_pp0_iter17_reg;
            do_cos_read_reg_1592_pp0_iter19_reg <= do_cos_read_reg_1592_pp0_iter18_reg;
            do_cos_read_reg_1592_pp0_iter20_reg <= do_cos_read_reg_1592_pp0_iter19_reg;
            do_cos_read_reg_1592_pp0_iter21_reg <= do_cos_read_reg_1592_pp0_iter20_reg;
            do_cos_read_reg_1592_pp0_iter22_reg <= do_cos_read_reg_1592_pp0_iter21_reg;
            do_cos_read_reg_1592_pp0_iter23_reg <= do_cos_read_reg_1592_pp0_iter22_reg;
            do_cos_read_reg_1592_pp0_iter24_reg <= do_cos_read_reg_1592_pp0_iter23_reg;
            do_cos_read_reg_1592_pp0_iter25_reg <= do_cos_read_reg_1592_pp0_iter24_reg;
            do_cos_read_reg_1592_pp0_iter26_reg <= do_cos_read_reg_1592_pp0_iter25_reg;
            do_cos_read_reg_1592_pp0_iter27_reg <= do_cos_read_reg_1592_pp0_iter26_reg;
            do_cos_read_reg_1592_pp0_iter28_reg <= do_cos_read_reg_1592_pp0_iter27_reg;
            do_cos_read_reg_1592_pp0_iter29_reg <= do_cos_read_reg_1592_pp0_iter28_reg;
            do_cos_read_reg_1592_pp0_iter2_reg <= do_cos_read_reg_1592_pp0_iter1_reg;
            do_cos_read_reg_1592_pp0_iter30_reg <= do_cos_read_reg_1592_pp0_iter29_reg;
            do_cos_read_reg_1592_pp0_iter3_reg <= do_cos_read_reg_1592_pp0_iter2_reg;
            do_cos_read_reg_1592_pp0_iter4_reg <= do_cos_read_reg_1592_pp0_iter3_reg;
            do_cos_read_reg_1592_pp0_iter5_reg <= do_cos_read_reg_1592_pp0_iter4_reg;
            do_cos_read_reg_1592_pp0_iter6_reg <= do_cos_read_reg_1592_pp0_iter5_reg;
            do_cos_read_reg_1592_pp0_iter7_reg <= do_cos_read_reg_1592_pp0_iter6_reg;
            do_cos_read_reg_1592_pp0_iter8_reg <= do_cos_read_reg_1592_pp0_iter7_reg;
            do_cos_read_reg_1592_pp0_iter9_reg <= do_cos_read_reg_1592_pp0_iter8_reg;
            fourth_order_double_sin_cos_K1_load_reg_1784 <= fourth_order_double_sin_cos_K1_q0;
            fourth_order_double_sin_cos_K2_load_reg_1789 <= fourth_order_double_sin_cos_K2_q0;
            fourth_order_double_sin_cos_K3_load_reg_1867 <= fourth_order_double_sin_cos_K3_q0;
            fourth_order_double_sin_cos_K4_load_reg_1877 <= fourth_order_double_sin_cos_K4_q0;
            h_reg_1657 <= grp_fu_380_p2;
            icmp_ln271_1_reg_1651 <= icmp_ln271_1_fu_479_p2;
            icmp_ln271_1_reg_1651_pp0_iter10_reg <= icmp_ln271_1_reg_1651_pp0_iter9_reg;
            icmp_ln271_1_reg_1651_pp0_iter11_reg <= icmp_ln271_1_reg_1651_pp0_iter10_reg;
            icmp_ln271_1_reg_1651_pp0_iter12_reg <= icmp_ln271_1_reg_1651_pp0_iter11_reg;
            icmp_ln271_1_reg_1651_pp0_iter13_reg <= icmp_ln271_1_reg_1651_pp0_iter12_reg;
            icmp_ln271_1_reg_1651_pp0_iter14_reg <= icmp_ln271_1_reg_1651_pp0_iter13_reg;
            icmp_ln271_1_reg_1651_pp0_iter15_reg <= icmp_ln271_1_reg_1651_pp0_iter14_reg;
            icmp_ln271_1_reg_1651_pp0_iter16_reg <= icmp_ln271_1_reg_1651_pp0_iter15_reg;
            icmp_ln271_1_reg_1651_pp0_iter17_reg <= icmp_ln271_1_reg_1651_pp0_iter16_reg;
            icmp_ln271_1_reg_1651_pp0_iter18_reg <= icmp_ln271_1_reg_1651_pp0_iter17_reg;
            icmp_ln271_1_reg_1651_pp0_iter19_reg <= icmp_ln271_1_reg_1651_pp0_iter18_reg;
            icmp_ln271_1_reg_1651_pp0_iter20_reg <= icmp_ln271_1_reg_1651_pp0_iter19_reg;
            icmp_ln271_1_reg_1651_pp0_iter21_reg <= icmp_ln271_1_reg_1651_pp0_iter20_reg;
            icmp_ln271_1_reg_1651_pp0_iter22_reg <= icmp_ln271_1_reg_1651_pp0_iter21_reg;
            icmp_ln271_1_reg_1651_pp0_iter23_reg <= icmp_ln271_1_reg_1651_pp0_iter22_reg;
            icmp_ln271_1_reg_1651_pp0_iter24_reg <= icmp_ln271_1_reg_1651_pp0_iter23_reg;
            icmp_ln271_1_reg_1651_pp0_iter25_reg <= icmp_ln271_1_reg_1651_pp0_iter24_reg;
            icmp_ln271_1_reg_1651_pp0_iter26_reg <= icmp_ln271_1_reg_1651_pp0_iter25_reg;
            icmp_ln271_1_reg_1651_pp0_iter27_reg <= icmp_ln271_1_reg_1651_pp0_iter26_reg;
            icmp_ln271_1_reg_1651_pp0_iter28_reg <= icmp_ln271_1_reg_1651_pp0_iter27_reg;
            icmp_ln271_1_reg_1651_pp0_iter29_reg <= icmp_ln271_1_reg_1651_pp0_iter28_reg;
            icmp_ln271_1_reg_1651_pp0_iter30_reg <= icmp_ln271_1_reg_1651_pp0_iter29_reg;
            icmp_ln271_1_reg_1651_pp0_iter31_reg <= icmp_ln271_1_reg_1651_pp0_iter30_reg;
            icmp_ln271_1_reg_1651_pp0_iter4_reg <= icmp_ln271_1_reg_1651;
            icmp_ln271_1_reg_1651_pp0_iter5_reg <= icmp_ln271_1_reg_1651_pp0_iter4_reg;
            icmp_ln271_1_reg_1651_pp0_iter6_reg <= icmp_ln271_1_reg_1651_pp0_iter5_reg;
            icmp_ln271_1_reg_1651_pp0_iter7_reg <= icmp_ln271_1_reg_1651_pp0_iter6_reg;
            icmp_ln271_1_reg_1651_pp0_iter8_reg <= icmp_ln271_1_reg_1651_pp0_iter7_reg;
            icmp_ln271_1_reg_1651_pp0_iter9_reg <= icmp_ln271_1_reg_1651_pp0_iter8_reg;
            icmp_ln271_reg_1714 <= icmp_ln271_fu_645_p2;
            icmp_ln271_reg_1714_pp0_iter10_reg <= icmp_ln271_reg_1714;
            icmp_ln271_reg_1714_pp0_iter11_reg <= icmp_ln271_reg_1714_pp0_iter10_reg;
            icmp_ln271_reg_1714_pp0_iter12_reg <= icmp_ln271_reg_1714_pp0_iter11_reg;
            icmp_ln271_reg_1714_pp0_iter13_reg <= icmp_ln271_reg_1714_pp0_iter12_reg;
            icmp_ln271_reg_1714_pp0_iter14_reg <= icmp_ln271_reg_1714_pp0_iter13_reg;
            icmp_ln271_reg_1714_pp0_iter15_reg <= icmp_ln271_reg_1714_pp0_iter14_reg;
            icmp_ln271_reg_1714_pp0_iter16_reg <= icmp_ln271_reg_1714_pp0_iter15_reg;
            icmp_ln271_reg_1714_pp0_iter17_reg <= icmp_ln271_reg_1714_pp0_iter16_reg;
            icmp_ln271_reg_1714_pp0_iter18_reg <= icmp_ln271_reg_1714_pp0_iter17_reg;
            icmp_ln271_reg_1714_pp0_iter19_reg <= icmp_ln271_reg_1714_pp0_iter18_reg;
            icmp_ln271_reg_1714_pp0_iter20_reg <= icmp_ln271_reg_1714_pp0_iter19_reg;
            icmp_ln271_reg_1714_pp0_iter21_reg <= icmp_ln271_reg_1714_pp0_iter20_reg;
            icmp_ln271_reg_1714_pp0_iter22_reg <= icmp_ln271_reg_1714_pp0_iter21_reg;
            icmp_ln271_reg_1714_pp0_iter23_reg <= icmp_ln271_reg_1714_pp0_iter22_reg;
            icmp_ln271_reg_1714_pp0_iter24_reg <= icmp_ln271_reg_1714_pp0_iter23_reg;
            icmp_ln271_reg_1714_pp0_iter25_reg <= icmp_ln271_reg_1714_pp0_iter24_reg;
            icmp_ln271_reg_1714_pp0_iter26_reg <= icmp_ln271_reg_1714_pp0_iter25_reg;
            icmp_ln271_reg_1714_pp0_iter27_reg <= icmp_ln271_reg_1714_pp0_iter26_reg;
            icmp_ln271_reg_1714_pp0_iter28_reg <= icmp_ln271_reg_1714_pp0_iter27_reg;
            icmp_ln271_reg_1714_pp0_iter29_reg <= icmp_ln271_reg_1714_pp0_iter28_reg;
            icmp_ln271_reg_1714_pp0_iter30_reg <= icmp_ln271_reg_1714_pp0_iter29_reg;
            icmp_ln271_reg_1714_pp0_iter31_reg <= icmp_ln271_reg_1714_pp0_iter30_reg;
            icmp_ln282_reg_1720 <= icmp_ln282_fu_650_p2;
            icmp_ln282_reg_1720_pp0_iter10_reg <= icmp_ln282_reg_1720;
            icmp_ln282_reg_1720_pp0_iter11_reg <= icmp_ln282_reg_1720_pp0_iter10_reg;
            icmp_ln282_reg_1720_pp0_iter12_reg <= icmp_ln282_reg_1720_pp0_iter11_reg;
            icmp_ln282_reg_1720_pp0_iter13_reg <= icmp_ln282_reg_1720_pp0_iter12_reg;
            icmp_ln282_reg_1720_pp0_iter14_reg <= icmp_ln282_reg_1720_pp0_iter13_reg;
            icmp_ln282_reg_1720_pp0_iter15_reg <= icmp_ln282_reg_1720_pp0_iter14_reg;
            icmp_ln282_reg_1720_pp0_iter16_reg <= icmp_ln282_reg_1720_pp0_iter15_reg;
            icmp_ln282_reg_1720_pp0_iter17_reg <= icmp_ln282_reg_1720_pp0_iter16_reg;
            icmp_ln282_reg_1720_pp0_iter18_reg <= icmp_ln282_reg_1720_pp0_iter17_reg;
            icmp_ln282_reg_1720_pp0_iter19_reg <= icmp_ln282_reg_1720_pp0_iter18_reg;
            icmp_ln282_reg_1720_pp0_iter20_reg <= icmp_ln282_reg_1720_pp0_iter19_reg;
            icmp_ln282_reg_1720_pp0_iter21_reg <= icmp_ln282_reg_1720_pp0_iter20_reg;
            icmp_ln282_reg_1720_pp0_iter22_reg <= icmp_ln282_reg_1720_pp0_iter21_reg;
            icmp_ln282_reg_1720_pp0_iter23_reg <= icmp_ln282_reg_1720_pp0_iter22_reg;
            icmp_ln282_reg_1720_pp0_iter24_reg <= icmp_ln282_reg_1720_pp0_iter23_reg;
            icmp_ln282_reg_1720_pp0_iter25_reg <= icmp_ln282_reg_1720_pp0_iter24_reg;
            icmp_ln282_reg_1720_pp0_iter26_reg <= icmp_ln282_reg_1720_pp0_iter25_reg;
            icmp_ln282_reg_1720_pp0_iter27_reg <= icmp_ln282_reg_1720_pp0_iter26_reg;
            icmp_ln282_reg_1720_pp0_iter28_reg <= icmp_ln282_reg_1720_pp0_iter27_reg;
            icmp_ln282_reg_1720_pp0_iter29_reg <= icmp_ln282_reg_1720_pp0_iter28_reg;
            icmp_ln282_reg_1720_pp0_iter30_reg <= icmp_ln282_reg_1720_pp0_iter29_reg;
            icmp_ln282_reg_1720_pp0_iter31_reg <= icmp_ln282_reg_1720_pp0_iter30_reg;
            icmp_ln424_1_reg_2004 <= icmp_ln424_1_fu_1299_p2;
            icmp_ln424_2_reg_2016 <= icmp_ln424_2_fu_1311_p2;
            icmp_ln424_reg_1985 <= icmp_ln424_fu_1279_p2;
            icmp_ln433_reg_1975 <= icmp_ln433_fu_1224_p2;
            icmp_ln433_reg_1975_pp0_iter30_reg <= icmp_ln433_reg_1975;
            in_shift_1_reg_1969 <= in_shift_1_fu_1219_p2;
            in_shift_1_reg_1969_pp0_iter30_reg <= in_shift_1_reg_1969;
            in_shift_2_reg_1998 <= in_shift_2_fu_1294_p2;
            in_shift_2_reg_1998_pp0_iter31_reg <= in_shift_2_reg_1998;
            in_shift_3_reg_2026 <= in_shift_3_fu_1355_p2;
            k_1_reg_1684 <= k_1_fu_598_p3;
            k_1_reg_1684_pp0_iter10_reg <= k_1_reg_1684;
            k_1_reg_1684_pp0_iter11_reg <= k_1_reg_1684_pp0_iter10_reg;
            k_1_reg_1684_pp0_iter12_reg <= k_1_reg_1684_pp0_iter11_reg;
            k_1_reg_1684_pp0_iter13_reg <= k_1_reg_1684_pp0_iter12_reg;
            k_reg_1668 <= {{grp_fu_380_p2[169:167]}};
            k_reg_1668_pp0_iter8_reg <= k_reg_1668;
            lshr_ln_reg_1907 <= {{grp_fu_348_p2[59:31]}};
            or_ln424_reg_2036 <= or_ln424_fu_1391_p2;
            or_ln433_reg_2041 <= or_ln433_fu_1434_p2;
            result_reg_1937 <= {{grp_fu_376_p2[125:63]}};
            results_exp_1_reg_2051 <= results_exp_1_fu_1496_p3;
            results_sign_3_reg_1773 <= results_sign_3_fu_945_p2;
            results_sign_4_reg_1800 <= results_sign_4_fu_975_p3;
            results_sign_4_reg_1800_pp0_iter16_reg <= results_sign_4_reg_1800;
            results_sign_4_reg_1800_pp0_iter17_reg <= results_sign_4_reg_1800_pp0_iter16_reg;
            results_sign_4_reg_1800_pp0_iter18_reg <= results_sign_4_reg_1800_pp0_iter17_reg;
            results_sign_4_reg_1800_pp0_iter19_reg <= results_sign_4_reg_1800_pp0_iter18_reg;
            results_sign_4_reg_1800_pp0_iter20_reg <= results_sign_4_reg_1800_pp0_iter19_reg;
            results_sign_4_reg_1800_pp0_iter21_reg <= results_sign_4_reg_1800_pp0_iter20_reg;
            results_sign_4_reg_1800_pp0_iter22_reg <= results_sign_4_reg_1800_pp0_iter21_reg;
            results_sign_4_reg_1800_pp0_iter23_reg <= results_sign_4_reg_1800_pp0_iter22_reg;
            results_sign_4_reg_1800_pp0_iter24_reg <= results_sign_4_reg_1800_pp0_iter23_reg;
            results_sign_4_reg_1800_pp0_iter25_reg <= results_sign_4_reg_1800_pp0_iter24_reg;
            results_sign_4_reg_1800_pp0_iter26_reg <= results_sign_4_reg_1800_pp0_iter25_reg;
            results_sign_4_reg_1800_pp0_iter27_reg <= results_sign_4_reg_1800_pp0_iter26_reg;
            results_sign_4_reg_1800_pp0_iter28_reg <= results_sign_4_reg_1800_pp0_iter27_reg;
            results_sign_4_reg_1800_pp0_iter29_reg <= results_sign_4_reg_1800_pp0_iter28_reg;
            results_sign_4_reg_1800_pp0_iter30_reg <= results_sign_4_reg_1800_pp0_iter29_reg;
            results_sign_4_reg_1800_pp0_iter31_reg <= results_sign_4_reg_1800_pp0_iter30_reg;
            select_ln424_4_reg_2046 <= select_ln424_4_fu_1458_p3;
            shift_1_reg_1993 <= shift_1_fu_1284_p2;
            shift_2_reg_2010 <= shift_2_fu_1305_p2;
            sub_ln506_reg_1709 <= sub_ln506_fu_639_p2;
            t1_reg_1847 <= fourth_order_double_sin_cos_K0_q0;
            tmp_10_reg_1862 <= {{grp_fu_364_p2[97:56]}};
            tmp_11_reg_1872 <= {{grp_fu_368_p2[97:63]}};
            tmp_12_reg_1912 <= {{grp_fu_352_p2[74:38]}};
            tmp_3_i_reg_1948 <= {{grp_fu_376_p2[109:94]}};
            tmp_3_i_reg_1948_pp0_iter29_reg <= tmp_3_i_reg_1948;
            tmp_3_reg_1703 <= Ex_1_fu_625_p2[32'd10];
            tmp_6_i_reg_1953 <= {{grp_fu_376_p2[93:78]}};
            tmp_6_i_reg_1953_pp0_iter29_reg <= tmp_6_i_reg_1953;
            tmp_8_reg_1728 <= {{x_1_fu_674_p3[62:56]}};
            tmp_8_reg_1728_pp0_iter11_reg <= tmp_8_reg_1728;
            tmp_8_reg_1728_pp0_iter12_reg <= tmp_8_reg_1728_pp0_iter11_reg;
            tmp_8_reg_1728_pp0_iter13_reg <= tmp_8_reg_1728_pp0_iter12_reg;
            tmp_9_i_reg_1958 <= {{grp_fu_376_p2[77:63]}};
            tmp_9_i_reg_1958_pp0_iter29_reg <= tmp_9_i_reg_1958;
            tmp_9_i_reg_1958_pp0_iter30_reg <= tmp_9_i_reg_1958_pp0_iter29_reg;
            tmp_i_reg_1943 <= {{grp_fu_376_p2[125:110]}};
            trunc_ln1_reg_1857 <= {{grp_fu_356_p2[92:45]}};
            trunc_ln_reg_1852 <= {{grp_fu_372_p2[107:52]}};
            zext_ln25_reg_1743[48 : 0] <= zext_ln25_fu_705_p1[48 : 0];
            zext_ln25_reg_1743_pp0_iter12_reg[48 : 0] <= zext_ln25_reg_1743[48 : 0];
            zext_ln25_reg_1743_pp0_iter13_reg[48 : 0] <= zext_ln25_reg_1743_pp0_iter12_reg[48 : 0];
            zext_ln25_reg_1743_pp0_iter14_reg[48 : 0] <= zext_ln25_reg_1743_pp0_iter13_reg[48 : 0];
            zext_ln25_reg_1743_pp0_iter15_reg[48 : 0] <= zext_ln25_reg_1743_pp0_iter14_reg[48 : 0];
            zext_ln32_reg_1756[7 : 0] <= zext_ln32_fu_776_p1[7 : 0];
            zext_ln32_reg_1756_pp0_iter15_reg[7 : 0] <= zext_ln32_reg_1756[7 : 0];
            zext_ln32_reg_1756_pp0_iter16_reg[7 : 0] <= zext_ln32_reg_1756_pp0_iter15_reg[7 : 0];
            zext_ln32_reg_1756_pp0_iter17_reg[7 : 0] <= zext_ln32_reg_1756_pp0_iter16_reg[7 : 0];
            zext_ln32_reg_1756_pp0_iter18_reg[7 : 0] <= zext_ln32_reg_1756_pp0_iter17_reg[7 : 0];
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            closepath_reg_1619 <= closepath_fu_410_p2;
            closepath_reg_1619_pp0_iter1_reg <= closepath_reg_1619;
            din_exp_reg_1606 <= {{data_fu_384_p1[62:52]}};
            din_exp_reg_1606_pp0_iter1_reg <= din_exp_reg_1606;
            din_sig_reg_1613 <= din_sig_fu_406_p1;
            din_sig_reg_1613_pp0_iter1_reg <= din_sig_reg_1613;
            din_sign_reg_1600 <= data_fu_384_p1[32'd63];
            din_sign_reg_1600_pp0_iter1_reg <= din_sign_reg_1600;
            do_cos_read_reg_1592 <= do_cos;
            do_cos_read_reg_1592_pp0_iter1_reg <= do_cos_read_reg_1592;
            table_256_reg_1636 <= ref_4oPi_table_256_q0;
            trunc_ln398_reg_1631 <= trunc_ln398_fu_445_p1;
            trunc_ln398_reg_1631_pp0_iter1_reg <= trunc_ln398_reg_1631;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter32 == 1'b1))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_idle_pp0 == 1'b1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter32 == 1'b0) 
    & (ap_enable_reg_pp0_iter31 == 1'b0) & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter26 == 1'b0) & (ap_enable_reg_pp0_iter25 == 1'b0) & (ap_enable_reg_pp0_iter24 == 1'b0) & (ap_enable_reg_pp0_iter23 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter31 == 1'b0) 
    & (ap_enable_reg_pp0_iter30 == 1'b0) & (ap_enable_reg_pp0_iter29 == 1'b0) & (ap_enable_reg_pp0_iter28 == 1'b0) & (ap_enable_reg_pp0_iter27 == 1'b0))) begin
            ap_idle_pp0_0to31 = 1'b1;
        end else begin
            ap_idle_pp0_0to31 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (ap_idle_pp0_0to31 == 1'b1))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            fourth_order_double_sin_cos_K0_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            fourth_order_double_sin_cos_K1_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter14 == 1'b1) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            fourth_order_double_sin_cos_K2_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            fourth_order_double_sin_cos_K3_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter19 == 1'b1) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            fourth_order_double_sin_cos_K4_ce0 = 1'b1;
        end else begin
            fourth_order_double_sin_cos_K4_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_348_ce = 1'b1;
        end else begin
            grp_fu_348_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_352_ce = 1'b1;
        end else begin
            grp_fu_352_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_356_ce = 1'b1;
        end else begin
            grp_fu_356_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_360_ce = 1'b1;
        end else begin
            grp_fu_360_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_364_ce = 1'b1;
        end else begin
            grp_fu_364_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_368_ce = 1'b1;
        end else begin
            grp_fu_368_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_372_ce = 1'b1;
        end else begin
            grp_fu_372_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_376_ce = 1'b1;
        end else begin
            grp_fu_376_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            grp_fu_380_ce = 1'b1;
        end else begin
            grp_fu_380_ce = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_ce) & (1'b0 == ap_block_pp0_stage0_11001))) begin
            ref_4oPi_table_256_ce0 = 1'b1;
        end else begin
            ref_4oPi_table_256_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign A_fu_769_p3 = {{sin_basis_fu_762_p3}, {tmp_8_reg_1728_pp0_iter13_reg}};

    assign B_fu_691_p1 = x_1_fu_674_p3[55:0];

    assign Ex_1_fu_625_p2 = (select_ln453_fu_591_p3 - zext_ln505_fu_604_p1);

    assign Ex_2_fu_1317_p3 = ((cos_basis_reg_1750_pp0_iter30_reg[0:0] == 1'b1) ? 11'd0 : Ex_1_reg_1697_pp0_iter30_reg);

    assign Ex_fu_586_p2 = ($signed(din_exp_reg_1606_pp0_iter8_reg) + $signed(11'd1027));

    assign Mx_1_fu_1109_p3 = ((cos_basis_reg_1750_pp0_iter22_reg[0:0] == 1'b1) ? 63'd9223372036854775807 : Mx_reg_1690_pp0_iter22_reg);

    assign Mx_bits_1_fu_522_p2 = (124'd0 - Mx_bits_reg_1662);

    assign Mx_bits_3_fu_527_p3 = ((and_ln451_fu_516_p2[0:0] == 1'b1) ? Mx_bits_1_fu_522_p2 : Mx_bits_reg_1662);

    assign Mx_zeros_fu_582_p1 = tmp_6_fu_574_p3[6:0];

    assign X_fu_467_p3 = {{1'd1}, {din_sig_reg_1613_pp0_iter2_reg}};

    assign add_ln37_1_fu_1083_p2 = ($signed(add_ln37_fu_1074_p2) + $signed(sext_ln37_2_fu_1080_p1));

    assign add_ln37_2_fu_1118_p2 = (add_ln37_1_reg_1902_pp0_iter22_reg + zext_ln37_2_fu_1115_p1);

    assign add_ln37_3_fu_1126_p2 = (add_ln37_2_fu_1118_p2 + zext_ln37_fu_1123_p1);

    assign add_ln37_fu_1074_p2 = ($signed(sext_ln37_fu_1067_p1) + $signed(sext_ln37_1_fu_1071_p1));

    assign add_ln396_fu_416_p2 = ($signed(din_exp_fu_396_p4) + $signed(11'd1101));

    assign add_ln422_fu_1360_p2 = (c_3_fu_1344_p3 + shift_2_reg_2010);

    assign add_ln432_fu_1410_p2 = ($signed(sext_ln252_fu_1323_p1) + $signed(12'd1023));

    assign addr_fu_422_p3 = ((closepath_fu_410_p2[0:0] == 1'b1) ? 11'd74 : add_ln396_fu_416_p2);

    assign and_ln271_1_fu_1550_p2 = (icmp_ln271_reg_1714_pp0_iter31_reg & icmp_ln271_1_reg_1651_pp0_iter31_reg);

    assign and_ln271_fu_961_p2 = (icmp_ln271_reg_1714_pp0_iter14_reg & icmp_ln271_1_reg_1651_pp0_iter14_reg);

    assign and_ln424_1_fu_1369_p2 = (icmp_ln424_reg_1985 & and_ln424_fu_1365_p2);

    assign and_ln424_2_fu_1379_p2 = (xor_ln424_fu_1374_p2 & icmp_ln424_reg_1985);

    assign and_ln424_fu_1365_p2 = (icmp_ln424_2_reg_2016 & icmp_ln424_1_reg_2004);

    assign and_ln451_fu_516_p2 = (xor_ln451_fu_511_p2 & tmp_fu_504_p3);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    always @(*) begin
        ap_block_pp0_stage0_subdone = (1'b0 == ap_ce);
    end

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_enable_reg_pp0_iter0 = ap_start;

    assign ap_return = t_2_fu_1580_p4;


    always @(tmp_5_i_fu_1243_p4) begin
        if (tmp_5_i_fu_1243_p4[0] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd0;
        end else if (tmp_5_i_fu_1243_p4[1] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd1;
        end else if (tmp_5_i_fu_1243_p4[2] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd2;
        end else if (tmp_5_i_fu_1243_p4[3] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd3;
        end else if (tmp_5_i_fu_1243_p4[4] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd4;
        end else if (tmp_5_i_fu_1243_p4[5] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd5;
        end else if (tmp_5_i_fu_1243_p4[6] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd6;
        end else if (tmp_5_i_fu_1243_p4[7] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd7;
        end else if (tmp_5_i_fu_1243_p4[8] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd8;
        end else if (tmp_5_i_fu_1243_p4[9] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd9;
        end else if (tmp_5_i_fu_1243_p4[10] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd10;
        end else if (tmp_5_i_fu_1243_p4[11] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd11;
        end else if (tmp_5_i_fu_1243_p4[12] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd12;
        end else if (tmp_5_i_fu_1243_p4[13] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd13;
        end else if (tmp_5_i_fu_1243_p4[14] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd14;
        end else if (tmp_5_i_fu_1243_p4[15] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd15;
        end else if (tmp_5_i_fu_1243_p4[16] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd16;
        end else if (tmp_5_i_fu_1243_p4[17] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd17;
        end else if (tmp_5_i_fu_1243_p4[18] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd18;
        end else if (tmp_5_i_fu_1243_p4[19] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd19;
        end else if (tmp_5_i_fu_1243_p4[20] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd20;
        end else if (tmp_5_i_fu_1243_p4[21] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd21;
        end else if (tmp_5_i_fu_1243_p4[22] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd22;
        end else if (tmp_5_i_fu_1243_p4[23] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd23;
        end else if (tmp_5_i_fu_1243_p4[24] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd24;
        end else if (tmp_5_i_fu_1243_p4[25] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd25;
        end else if (tmp_5_i_fu_1243_p4[26] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd26;
        end else if (tmp_5_i_fu_1243_p4[27] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd27;
        end else if (tmp_5_i_fu_1243_p4[28] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd28;
        end else if (tmp_5_i_fu_1243_p4[29] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd29;
        end else if (tmp_5_i_fu_1243_p4[30] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd30;
        end else if (tmp_5_i_fu_1243_p4[31] == 1'b1) begin
            c_1_fu_1253_p3 = 32'd31;
        end else begin
            c_1_fu_1253_p3 = 32'd32;
        end
    end


    always @(tmp_8_i_fu_1261_p4) begin
        if (tmp_8_i_fu_1261_p4[0] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd0;
        end else if (tmp_8_i_fu_1261_p4[1] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd1;
        end else if (tmp_8_i_fu_1261_p4[2] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd2;
        end else if (tmp_8_i_fu_1261_p4[3] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd3;
        end else if (tmp_8_i_fu_1261_p4[4] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd4;
        end else if (tmp_8_i_fu_1261_p4[5] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd5;
        end else if (tmp_8_i_fu_1261_p4[6] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd6;
        end else if (tmp_8_i_fu_1261_p4[7] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd7;
        end else if (tmp_8_i_fu_1261_p4[8] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd8;
        end else if (tmp_8_i_fu_1261_p4[9] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd9;
        end else if (tmp_8_i_fu_1261_p4[10] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd10;
        end else if (tmp_8_i_fu_1261_p4[11] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd11;
        end else if (tmp_8_i_fu_1261_p4[12] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd12;
        end else if (tmp_8_i_fu_1261_p4[13] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd13;
        end else if (tmp_8_i_fu_1261_p4[14] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd14;
        end else if (tmp_8_i_fu_1261_p4[15] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd15;
        end else if (tmp_8_i_fu_1261_p4[16] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd16;
        end else if (tmp_8_i_fu_1261_p4[17] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd17;
        end else if (tmp_8_i_fu_1261_p4[18] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd18;
        end else if (tmp_8_i_fu_1261_p4[19] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd19;
        end else if (tmp_8_i_fu_1261_p4[20] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd20;
        end else if (tmp_8_i_fu_1261_p4[21] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd21;
        end else if (tmp_8_i_fu_1261_p4[22] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd22;
        end else if (tmp_8_i_fu_1261_p4[23] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd23;
        end else if (tmp_8_i_fu_1261_p4[24] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd24;
        end else if (tmp_8_i_fu_1261_p4[25] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd25;
        end else if (tmp_8_i_fu_1261_p4[26] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd26;
        end else if (tmp_8_i_fu_1261_p4[27] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd27;
        end else if (tmp_8_i_fu_1261_p4[28] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd28;
        end else if (tmp_8_i_fu_1261_p4[29] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd29;
        end else if (tmp_8_i_fu_1261_p4[30] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd30;
        end else if (tmp_8_i_fu_1261_p4[31] == 1'b1) begin
            c_2_fu_1271_p3 = 32'd31;
        end else begin
            c_2_fu_1271_p3 = 32'd32;
        end
    end


    always @(tmp_i_63_fu_1334_p4) begin
        if (tmp_i_63_fu_1334_p4[0] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd0;
        end else if (tmp_i_63_fu_1334_p4[1] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd1;
        end else if (tmp_i_63_fu_1334_p4[2] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd2;
        end else if (tmp_i_63_fu_1334_p4[3] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd3;
        end else if (tmp_i_63_fu_1334_p4[4] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd4;
        end else if (tmp_i_63_fu_1334_p4[5] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd5;
        end else if (tmp_i_63_fu_1334_p4[6] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd6;
        end else if (tmp_i_63_fu_1334_p4[7] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd7;
        end else if (tmp_i_63_fu_1334_p4[8] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd8;
        end else if (tmp_i_63_fu_1334_p4[9] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd9;
        end else if (tmp_i_63_fu_1334_p4[10] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd10;
        end else if (tmp_i_63_fu_1334_p4[11] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd11;
        end else if (tmp_i_63_fu_1334_p4[12] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd12;
        end else if (tmp_i_63_fu_1334_p4[13] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd13;
        end else if (tmp_i_63_fu_1334_p4[14] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd14;
        end else if (tmp_i_63_fu_1334_p4[15] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd15;
        end else if (tmp_i_63_fu_1334_p4[16] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd16;
        end else if (tmp_i_63_fu_1334_p4[17] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd17;
        end else if (tmp_i_63_fu_1334_p4[18] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd18;
        end else if (tmp_i_63_fu_1334_p4[19] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd19;
        end else if (tmp_i_63_fu_1334_p4[20] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd20;
        end else if (tmp_i_63_fu_1334_p4[21] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd21;
        end else if (tmp_i_63_fu_1334_p4[22] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd22;
        end else if (tmp_i_63_fu_1334_p4[23] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd23;
        end else if (tmp_i_63_fu_1334_p4[24] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd24;
        end else if (tmp_i_63_fu_1334_p4[25] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd25;
        end else if (tmp_i_63_fu_1334_p4[26] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd26;
        end else if (tmp_i_63_fu_1334_p4[27] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd27;
        end else if (tmp_i_63_fu_1334_p4[28] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd28;
        end else if (tmp_i_63_fu_1334_p4[29] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd29;
        end else if (tmp_i_63_fu_1334_p4[30] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd30;
        end else if (tmp_i_63_fu_1334_p4[31] == 1'b1) begin
            c_3_fu_1344_p3 = 32'd31;
        end else begin
            c_3_fu_1344_p3 = 32'd32;
        end
    end


    always @(tmp_2_i_fu_1197_p4) begin
        if (tmp_2_i_fu_1197_p4[0] == 1'b1) begin
            c_fu_1207_p3 = 32'd0;
        end else if (tmp_2_i_fu_1197_p4[1] == 1'b1) begin
            c_fu_1207_p3 = 32'd1;
        end else if (tmp_2_i_fu_1197_p4[2] == 1'b1) begin
            c_fu_1207_p3 = 32'd2;
        end else if (tmp_2_i_fu_1197_p4[3] == 1'b1) begin
            c_fu_1207_p3 = 32'd3;
        end else if (tmp_2_i_fu_1197_p4[4] == 1'b1) begin
            c_fu_1207_p3 = 32'd4;
        end else if (tmp_2_i_fu_1197_p4[5] == 1'b1) begin
            c_fu_1207_p3 = 32'd5;
        end else if (tmp_2_i_fu_1197_p4[6] == 1'b1) begin
            c_fu_1207_p3 = 32'd6;
        end else if (tmp_2_i_fu_1197_p4[7] == 1'b1) begin
            c_fu_1207_p3 = 32'd7;
        end else if (tmp_2_i_fu_1197_p4[8] == 1'b1) begin
            c_fu_1207_p3 = 32'd8;
        end else if (tmp_2_i_fu_1197_p4[9] == 1'b1) begin
            c_fu_1207_p3 = 32'd9;
        end else if (tmp_2_i_fu_1197_p4[10] == 1'b1) begin
            c_fu_1207_p3 = 32'd10;
        end else if (tmp_2_i_fu_1197_p4[11] == 1'b1) begin
            c_fu_1207_p3 = 32'd11;
        end else if (tmp_2_i_fu_1197_p4[12] == 1'b1) begin
            c_fu_1207_p3 = 32'd12;
        end else if (tmp_2_i_fu_1197_p4[13] == 1'b1) begin
            c_fu_1207_p3 = 32'd13;
        end else if (tmp_2_i_fu_1197_p4[14] == 1'b1) begin
            c_fu_1207_p3 = 32'd14;
        end else if (tmp_2_i_fu_1197_p4[15] == 1'b1) begin
            c_fu_1207_p3 = 32'd15;
        end else if (tmp_2_i_fu_1197_p4[16] == 1'b1) begin
            c_fu_1207_p3 = 32'd16;
        end else if (tmp_2_i_fu_1197_p4[17] == 1'b1) begin
            c_fu_1207_p3 = 32'd17;
        end else if (tmp_2_i_fu_1197_p4[18] == 1'b1) begin
            c_fu_1207_p3 = 32'd18;
        end else if (tmp_2_i_fu_1197_p4[19] == 1'b1) begin
            c_fu_1207_p3 = 32'd19;
        end else if (tmp_2_i_fu_1197_p4[20] == 1'b1) begin
            c_fu_1207_p3 = 32'd20;
        end else if (tmp_2_i_fu_1197_p4[21] == 1'b1) begin
            c_fu_1207_p3 = 32'd21;
        end else if (tmp_2_i_fu_1197_p4[22] == 1'b1) begin
            c_fu_1207_p3 = 32'd22;
        end else if (tmp_2_i_fu_1197_p4[23] == 1'b1) begin
            c_fu_1207_p3 = 32'd23;
        end else if (tmp_2_i_fu_1197_p4[24] == 1'b1) begin
            c_fu_1207_p3 = 32'd24;
        end else if (tmp_2_i_fu_1197_p4[25] == 1'b1) begin
            c_fu_1207_p3 = 32'd25;
        end else if (tmp_2_i_fu_1197_p4[26] == 1'b1) begin
            c_fu_1207_p3 = 32'd26;
        end else if (tmp_2_i_fu_1197_p4[27] == 1'b1) begin
            c_fu_1207_p3 = 32'd27;
        end else if (tmp_2_i_fu_1197_p4[28] == 1'b1) begin
            c_fu_1207_p3 = 32'd28;
        end else if (tmp_2_i_fu_1197_p4[29] == 1'b1) begin
            c_fu_1207_p3 = 32'd29;
        end else if (tmp_2_i_fu_1197_p4[30] == 1'b1) begin
            c_fu_1207_p3 = 32'd30;
        end else if (tmp_2_i_fu_1197_p4[31] == 1'b1) begin
            c_fu_1207_p3 = 32'd31;
        end else begin
            c_fu_1207_p3 = 32'd32;
        end
    end

    assign closepath_fu_410_p2 = ((din_exp_fu_396_p4 < 11'd1022) ? 1'b1 : 1'b0);

    assign cos_basis_fu_755_p3 = ((do_cos_read_reg_1592_pp0_iter13_reg[0:0] == 1'b1) ? xor_ln242_fu_749_p2 : tmp_7_fu_710_p19);

    assign data_fu_384_p1 = t_in;

    assign din_exp_fu_396_p4 = {{data_fu_384_p1[62:52]}};

    assign din_sig_fu_406_p1 = data_fu_384_p1[51:0];

    assign empty_fu_1465_p1 = newexp_fu_1420_p2[10:0];

    assign fourth_order_double_sin_cos_K0_address0 = zext_ln32_reg_1756_pp0_iter18_reg;

    assign fourth_order_double_sin_cos_K1_address0 = zext_ln32_fu_776_p1;

    assign fourth_order_double_sin_cos_K2_address0 = zext_ln32_fu_776_p1;

    assign fourth_order_double_sin_cos_K3_address0 = zext_ln32_reg_1756_pp0_iter18_reg;

    assign fourth_order_double_sin_cos_K4_address0 = zext_ln32_reg_1756_pp0_iter18_reg;

    assign grp_fu_348_p0 = grp_fu_348_p00;

    assign grp_fu_348_p00 = tmp_11_reg_1872;

    assign grp_fu_348_p1 = grp_fu_348_p10;

    assign grp_fu_348_p10 = fourth_order_double_sin_cos_K4_load_reg_1877;

    assign grp_fu_352_p0 = grp_fu_352_p00;

    assign grp_fu_352_p00 = tmp_10_reg_1862;

    assign grp_fu_352_p1 = grp_fu_352_p10;

    assign grp_fu_352_p10 = fourth_order_double_sin_cos_K3_load_reg_1867;

    assign grp_fu_356_p0 = grp_fu_356_p00;

    assign grp_fu_356_p00 = B_squared_reg_1778;

    assign grp_fu_360_p0 = zext_ln25_fu_705_p1;

    assign grp_fu_360_p1 = zext_ln25_fu_705_p1;

    assign grp_fu_364_p0 = zext_ln25_1_fu_982_p1;

    assign grp_fu_364_p1 = zext_ln25_reg_1743_pp0_iter15_reg;

    assign grp_fu_368_p0 = zext_ln25_1_fu_982_p1;

    assign grp_fu_368_p1 = zext_ln25_1_fu_982_p1;

    assign grp_fu_372_p0 = grp_fu_372_p00;

    assign grp_fu_372_p00 = B_reg_1733_pp0_iter15_reg;

    assign grp_fu_376_p1 = grp_fu_376_p10;

    assign grp_fu_376_p10 = Mx_1_reg_1917;

    assign grp_fu_380_p1 = grp_fu_380_p10;

    assign grp_fu_380_p10 = X_fu_467_p3;

    assign icmp_ln271_1_fu_479_p2 = ((din_sig_reg_1613_pp0_iter2_reg == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln271_fu_645_p2 = ((din_exp_reg_1606_pp0_iter8_reg == 11'd0) ? 1'b1 : 1'b0);

    assign icmp_ln282_fu_650_p2 = ((din_exp_reg_1606_pp0_iter8_reg == 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln424_1_fu_1299_p2 = ((c_1_fu_1253_p3 == 32'd16) ? 1'b1 : 1'b0);

    assign icmp_ln424_2_fu_1311_p2 = ((c_2_fu_1271_p3 == 32'd16) ? 1'b1 : 1'b0);

    assign icmp_ln424_fu_1279_p2 = ((c_reg_1963 == 32'd16) ? 1'b1 : 1'b0);

    assign icmp_ln433_fu_1224_p2 = ((result_reg_1937 == 63'd0) ? 1'b1 : 1'b0);

    assign in_shift_1_fu_1219_p2 = result_reg_1937 << zext_ln423_fu_1215_p1;

    assign in_shift_2_fu_1294_p2 = in_shift_1_reg_1969 << zext_ln423_1_fu_1290_p1;

    assign in_shift_3_fu_1355_p2 = in_shift_2_reg_1998 << zext_ln423_2_fu_1352_p1;

    assign index_fu_782_p3 = {{din_sign_reg_1600_pp0_iter13_reg}, {k_1_reg_1684_pp0_iter13_reg}};

    assign k_1_fu_598_p3 = ((closepath_reg_1619_pp0_iter8_reg[0:0] == 1'b1) ? 3'd0 : k_reg_1668_pp0_iter8_reg);

    assign lshr_ln506_fu_664_p2 = Mx_reg_1690 >> zext_ln506_fu_660_p1;

    assign newexp_fu_1420_p2 = ($signed(
        sext_ln432_fu_1416_p1
    ) - $signed(
        select_ln424_2_fu_1402_p3
    ));

    assign or_ln271_fu_1568_p2 = (icmp_ln282_reg_1720_pp0_iter31_reg | and_ln271_reg_1794_pp0_iter31_reg);

    assign or_ln282_fu_1483_p2 = (or_ln433_fu_1434_p2 | icmp_ln282_reg_1720_pp0_iter30_reg);

    assign or_ln424_fu_1391_p2 = (and_ln424_2_fu_1379_p2 | and_ln424_1_fu_1369_p2);

    assign or_ln433_fu_1434_p2 = (tmp_13_fu_1426_p3 | icmp_ln433_reg_1975_pp0_iter30_reg);

    assign out_bits_4_fu_1229_p3 = {{tmp_3_i_reg_1948_pp0_iter29_reg}, {16'd32768}};

    assign out_bits_5_fu_1236_p3 = {{tmp_6_i_reg_1953_pp0_iter29_reg}, {16'd32768}};

    assign out_bits_6_fu_1327_p3 = {{tmp_9_i_reg_1958_pp0_iter30_reg}, {17'd65536}};

    assign out_bits_fu_1190_p3 = {{tmp_i_reg_1943}, {16'd32768}};

    assign ref_4oPi_table_256_address0 = zext_ln397_fu_440_p1;

    assign results_exp_1_fu_1496_p3 = ((and_ln271_reg_1794_pp0_iter30_reg[0:0] == 1'b1) ? select_ln259_fu_1469_p3 : results_exp_fu_1488_p3);

    assign results_exp_fu_1488_p3 = ((or_ln282_fu_1483_p2[0:0] == 1'b1) ? select_ln282_fu_1476_p3 : empty_fu_1465_p1);

    assign results_sig_1_fu_1572_p3 = ((or_ln271_fu_1568_p2[0:0] == 1'b1) ? select_ln271_fu_1560_p3 : significand_fu_1543_p3);

    assign results_sign_2_fu_970_p2 = (xor_ln278_fu_965_p2 & din_sign_reg_1600_pp0_iter14_reg);

    assign results_sign_3_fu_945_p2 = (xor_ln282_fu_940_p2 & results_sign_fu_932_p3);

    assign results_sign_4_fu_975_p3 = ((and_ln271_fu_961_p2[0:0] == 1'b1) ? results_sign_2_fu_970_p2 : results_sign_3_reg_1773);

    assign results_sign_fu_932_p3 = ((cos_basis_fu_755_p3[0:0] == 1'b1) ? tmp_9_fu_788_p35 : tmp_2_fu_860_p35);

    assign select_ln259_fu_1469_p3 = ((do_cos_read_reg_1592_pp0_iter30_reg[0:0] == 1'b1) ? 11'd1023 : 11'd0);

    assign select_ln271_fu_1560_p3 = ((xor_ln271_fu_1554_p2[0:0] == 1'b1) ? 52'd4503599627370495 : 52'd0);

    assign select_ln282_fu_1476_p3 = ((icmp_ln282_reg_1720_pp0_iter30_reg[0:0] == 1'b1) ? 11'd2047 : 11'd0);

    assign select_ln424_1_fu_1397_p3 = ((icmp_ln424_reg_1985[0:0] == 1'b1) ? shift_2_reg_2010 : c_reg_1963_pp0_iter30_reg);

    assign select_ln424_2_fu_1402_p3 = ((or_ln424_fu_1391_p2[0:0] == 1'b1) ? select_ln424_fu_1384_p3 : select_ln424_1_fu_1397_p3);

    assign select_ln424_3_fu_1530_p3 = ((and_ln424_2_reg_2031[0:0] == 1'b1) ? tmp_14_fu_1511_p4 : tmp_15_fu_1520_p4);

    assign select_ln424_4_fu_1458_p3 = ((icmp_ln424_reg_1985[0:0] == 1'b1) ? tmp_16_fu_1439_p4 : tmp_17_fu_1449_p4);

    assign select_ln424_5_fu_1537_p3 = ((or_ln424_reg_2036[0:0] == 1'b1) ? select_ln424_3_fu_1530_p3 : select_ln424_4_reg_2046);

    assign select_ln424_fu_1384_p3 = ((and_ln424_2_fu_1379_p2[0:0] == 1'b1) ? shift_1_reg_1993 : add_ln422_fu_1360_p2);

    assign select_ln453_fu_591_p3 = ((closepath_reg_1619_pp0_iter8_reg[0:0] == 1'b1) ? Ex_fu_586_p2 : 11'd0);

    assign select_ln506_fu_655_p3 = ((tmp_3_reg_1703[0:0] == 1'b1) ? sub_ln506_reg_1709 : Ex_1_reg_1697);

    assign sext_ln252_fu_1323_p1 = $signed(Ex_2_fu_1317_p3);

    assign sext_ln37_1_fu_1071_p1 = $signed(trunc_ln_reg_1852);

    assign sext_ln37_2_fu_1080_p1 = $signed(trunc_ln1_reg_1857);

    assign sext_ln37_fu_1067_p1 = $signed(t1_1_fu_1044_p3);

    assign sext_ln432_fu_1416_p1 = $signed(add_ln432_fu_1410_p2);

    assign sext_ln75_fu_570_p1 = $signed(tmp_5_fu_562_p3);

    assign shift_1_fu_1284_p2 = (c_1_fu_1253_p3 + 32'd16);

    assign shift_2_fu_1305_p2 = (c_2_fu_1271_p3 + shift_1_fu_1284_p2);

    assign shl_ln398_fu_452_p2 = table_256_reg_1636 << zext_ln398_fu_449_p1;

    assign shl_ln423_fu_1506_p2 = in_shift_3_reg_2026 << zext_ln423_3_fu_1503_p1;

    assign shl_ln504_fu_610_p2 = Mx_bits_3_reg_1673 << zext_ln504_fu_607_p1;

    assign shl_ln506_fu_669_p2 = Mx_reg_1690 << zext_ln506_fu_660_p1;

    assign significand_fu_1543_p3 = ((or_ln433_reg_2041[0:0] == 1'b1) ? 52'd0 : select_ln424_5_fu_1537_p3);

    assign sin_basis_fu_762_p3 = ((do_cos_read_reg_1592_pp0_iter13_reg[0:0] == 1'b1) ? tmp_7_fu_710_p19 : xor_ln242_fu_749_p2);

    assign sub_ln506_fu_639_p2 = (11'd0 - Ex_1_fu_625_p2);

    assign t1_1_fu_1044_p3 = {{t1_reg_1847}, {4'd0}};

    assign t_2_fu_1580_p4 = {
        {{results_sign_4_reg_1800_pp0_iter31_reg}, {results_exp_1_reg_2051}},
        {results_sig_1_fu_1572_p3}
    };

    assign t_fu_544_p3 = {{tmp_1_fu_534_p4}, {1'd1}};

    assign tmp_13_fu_1426_p3 = newexp_fu_1420_p2[32'd31];

    assign tmp_14_fu_1511_p4 = {{in_shift_2_reg_1998_pp0_iter31_reg[61:10]}};

    assign tmp_15_fu_1520_p4 = {{shl_ln423_fu_1506_p2[61:10]}};

    assign tmp_16_fu_1439_p4 = {{in_shift_3_fu_1355_p2[61:10]}};

    assign tmp_17_fu_1449_p4 = {{in_shift_1_reg_1969_pp0_iter30_reg[61:10]}};

    assign tmp_1_fu_534_p4 = {{Mx_bits_3_fu_527_p3[123:63]}};

    assign tmp_2_fu_860_p33 = 'bx;

    integer ap_tvar_int_0;

    always @(out_bits_fu_1190_p3) begin
        for (ap_tvar_int_0 = 32 - 1; ap_tvar_int_0 >= 0; ap_tvar_int_0 = ap_tvar_int_0 - 1) begin
            if (ap_tvar_int_0 > 31 - 0) begin
                tmp_2_i_fu_1197_p4[ap_tvar_int_0] = 1'b0;
            end else begin
                tmp_2_i_fu_1197_p4[ap_tvar_int_0] = out_bits_fu_1190_p3[31-ap_tvar_int_0];
            end
        end
    end

    integer ap_tvar_int_1;

    always @(t_fu_544_p3) begin
        for (ap_tvar_int_1 = 62 - 1; ap_tvar_int_1 >= 0; ap_tvar_int_1 = ap_tvar_int_1 - 1) begin
            if (ap_tvar_int_1 > 61 - 0) begin
                tmp_4_fu_552_p4[ap_tvar_int_1] = 1'b0;
            end else begin
                tmp_4_fu_552_p4[ap_tvar_int_1] = t_fu_544_p3[61-ap_tvar_int_1];
            end
        end
    end

    assign tmp_5_fu_562_p3 = {{1'd1}, {tmp_4_fu_552_p4}};

    integer ap_tvar_int_2;

    always @(out_bits_4_fu_1229_p3) begin
        for (ap_tvar_int_2 = 32 - 1; ap_tvar_int_2 >= 0; ap_tvar_int_2 = ap_tvar_int_2 - 1) begin
            if (ap_tvar_int_2 > 31 - 0) begin
                tmp_5_i_fu_1243_p4[ap_tvar_int_2] = 1'b0;
            end else begin
                tmp_5_i_fu_1243_p4[ap_tvar_int_2] = out_bits_4_fu_1229_p3[31-ap_tvar_int_2];
            end
        end
    end


    always @(sext_ln75_fu_570_p1) begin
        if (sext_ln75_fu_570_p1[0] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd0;
        end else if (sext_ln75_fu_570_p1[1] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd1;
        end else if (sext_ln75_fu_570_p1[2] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd2;
        end else if (sext_ln75_fu_570_p1[3] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd3;
        end else if (sext_ln75_fu_570_p1[4] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd4;
        end else if (sext_ln75_fu_570_p1[5] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd5;
        end else if (sext_ln75_fu_570_p1[6] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd6;
        end else if (sext_ln75_fu_570_p1[7] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd7;
        end else if (sext_ln75_fu_570_p1[8] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd8;
        end else if (sext_ln75_fu_570_p1[9] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd9;
        end else if (sext_ln75_fu_570_p1[10] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd10;
        end else if (sext_ln75_fu_570_p1[11] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd11;
        end else if (sext_ln75_fu_570_p1[12] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd12;
        end else if (sext_ln75_fu_570_p1[13] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd13;
        end else if (sext_ln75_fu_570_p1[14] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd14;
        end else if (sext_ln75_fu_570_p1[15] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd15;
        end else if (sext_ln75_fu_570_p1[16] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd16;
        end else if (sext_ln75_fu_570_p1[17] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd17;
        end else if (sext_ln75_fu_570_p1[18] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd18;
        end else if (sext_ln75_fu_570_p1[19] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd19;
        end else if (sext_ln75_fu_570_p1[20] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd20;
        end else if (sext_ln75_fu_570_p1[21] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd21;
        end else if (sext_ln75_fu_570_p1[22] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd22;
        end else if (sext_ln75_fu_570_p1[23] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd23;
        end else if (sext_ln75_fu_570_p1[24] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd24;
        end else if (sext_ln75_fu_570_p1[25] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd25;
        end else if (sext_ln75_fu_570_p1[26] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd26;
        end else if (sext_ln75_fu_570_p1[27] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd27;
        end else if (sext_ln75_fu_570_p1[28] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd28;
        end else if (sext_ln75_fu_570_p1[29] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd29;
        end else if (sext_ln75_fu_570_p1[30] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd30;
        end else if (sext_ln75_fu_570_p1[31] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd31;
        end else if (sext_ln75_fu_570_p1[32] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd32;
        end else if (sext_ln75_fu_570_p1[33] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd33;
        end else if (sext_ln75_fu_570_p1[34] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd34;
        end else if (sext_ln75_fu_570_p1[35] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd35;
        end else if (sext_ln75_fu_570_p1[36] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd36;
        end else if (sext_ln75_fu_570_p1[37] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd37;
        end else if (sext_ln75_fu_570_p1[38] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd38;
        end else if (sext_ln75_fu_570_p1[39] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd39;
        end else if (sext_ln75_fu_570_p1[40] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd40;
        end else if (sext_ln75_fu_570_p1[41] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd41;
        end else if (sext_ln75_fu_570_p1[42] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd42;
        end else if (sext_ln75_fu_570_p1[43] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd43;
        end else if (sext_ln75_fu_570_p1[44] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd44;
        end else if (sext_ln75_fu_570_p1[45] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd45;
        end else if (sext_ln75_fu_570_p1[46] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd46;
        end else if (sext_ln75_fu_570_p1[47] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd47;
        end else if (sext_ln75_fu_570_p1[48] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd48;
        end else if (sext_ln75_fu_570_p1[49] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd49;
        end else if (sext_ln75_fu_570_p1[50] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd50;
        end else if (sext_ln75_fu_570_p1[51] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd51;
        end else if (sext_ln75_fu_570_p1[52] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd52;
        end else if (sext_ln75_fu_570_p1[53] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd53;
        end else if (sext_ln75_fu_570_p1[54] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd54;
        end else if (sext_ln75_fu_570_p1[55] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd55;
        end else if (sext_ln75_fu_570_p1[56] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd56;
        end else if (sext_ln75_fu_570_p1[57] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd57;
        end else if (sext_ln75_fu_570_p1[58] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd58;
        end else if (sext_ln75_fu_570_p1[59] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd59;
        end else if (sext_ln75_fu_570_p1[60] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd60;
        end else if (sext_ln75_fu_570_p1[61] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd61;
        end else if (sext_ln75_fu_570_p1[62] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd62;
        end else if (sext_ln75_fu_570_p1[63] == 1'b1) begin
            tmp_6_fu_574_p3 = 64'd63;
        end else begin
            tmp_6_fu_574_p3 = 64'd64;
        end
    end

    assign tmp_7_fu_710_p17 = 'bx;

    integer ap_tvar_int_3;

    always @(out_bits_5_fu_1236_p3) begin
        for (ap_tvar_int_3 = 32 - 1; ap_tvar_int_3 >= 0; ap_tvar_int_3 = ap_tvar_int_3 - 1) begin
            if (ap_tvar_int_3 > 31 - 0) begin
                tmp_8_i_fu_1261_p4[ap_tvar_int_3] = 1'b0;
            end else begin
                tmp_8_i_fu_1261_p4[ap_tvar_int_3] = out_bits_5_fu_1236_p3[31-ap_tvar_int_3];
            end
        end
    end

    assign tmp_9_fu_788_p33 = 'bx;

    assign tmp_fu_504_p3 = h_reg_1657[32'd167];

    integer ap_tvar_int_4;

    always @(out_bits_6_fu_1327_p3) begin
        for (ap_tvar_int_4 = 32 - 1; ap_tvar_int_4 >= 0; ap_tvar_int_4 = ap_tvar_int_4 - 1) begin
            if (ap_tvar_int_4 > 31 - 0) begin
                tmp_i_63_fu_1334_p4[ap_tvar_int_4] = 1'b0;
            end else begin
                tmp_i_63_fu_1334_p4[ap_tvar_int_4] = out_bits_6_fu_1327_p3[31-ap_tvar_int_4];
            end
        end
    end

    assign tmp_s_fu_430_p4 = {{addr_fu_422_p3[10:7]}};

    assign trunc_ln398_fu_445_p1 = addr_fu_422_p3[6:0];

    assign x_1_fu_674_p3 = ((tmp_3_reg_1703[0:0] == 1'b1) ? lshr_ln506_fu_664_p2 : shl_ln506_fu_669_p2);

    assign xor_ln242_fu_749_p2 = (tmp_7_fu_710_p19 ^ 1'd1);

    assign xor_ln271_fu_1554_p2 = (1'd1 ^ and_ln271_1_fu_1550_p2);

    assign xor_ln278_fu_965_p2 = (do_cos_read_reg_1592_pp0_iter14_reg ^ 1'd1);

    assign xor_ln282_fu_940_p2 = (icmp_ln282_reg_1720_pp0_iter13_reg ^ 1'd1);

    assign xor_ln424_fu_1374_p2 = (icmp_ln424_1_reg_2004 ^ 1'd1);

    assign xor_ln451_fu_511_p2 = (closepath_reg_1619_pp0_iter7_reg ^ 1'd1);

    assign zext_ln25_1_fu_982_p1 = B_squared_reg_1778;

    assign zext_ln25_fu_705_p1 = B_trunc_reg_1738;

    assign zext_ln32_fu_776_p1 = A_fu_769_p3;

    assign zext_ln37_2_fu_1115_p1 = tmp_12_reg_1912;

    assign zext_ln37_fu_1123_p1 = lshr_ln_reg_1907;

    assign zext_ln397_fu_440_p1 = tmp_s_fu_430_p4;

    assign zext_ln398_fu_449_p1 = trunc_ln398_reg_1631_pp0_iter1_reg;

    assign zext_ln423_1_fu_1290_p1 = c_1_fu_1253_p3;

    assign zext_ln423_2_fu_1352_p1 = c_2_reg_1980;

    assign zext_ln423_3_fu_1503_p1 = c_3_reg_2021;

    assign zext_ln423_fu_1215_p1 = c_fu_1207_p3;

    assign zext_ln504_fu_607_p1 = Mx_zeros_reg_1678;

    assign zext_ln505_fu_604_p1 = Mx_zeros_reg_1678;

    assign zext_ln506_fu_660_p1 = select_ln506_fu_655_p3;

    always @(posedge ap_clk) begin
        zext_ln25_reg_1743[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln25_reg_1743_pp0_iter12_reg[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln25_reg_1743_pp0_iter13_reg[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln25_reg_1743_pp0_iter14_reg[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln25_reg_1743_pp0_iter15_reg[97:49] <= 49'b0000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1756[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1756_pp0_iter15_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1756_pp0_iter16_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1756_pp0_iter17_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
        zext_ln32_reg_1756_pp0_iter18_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    end

endmodule  //main_sin_or_cos_double_s
