/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1 (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    minDist,
    sub_ln296,
    rrtVertices_address0,
    rrtVertices_ce0,
    rrtVertices_q0,
    qRand_address0,
    qRand_ce0,
    qRand_q0,
    bestIdx_3_out,
    bestIdx_3_out_ap_vld,
    grp_fu_2529_p_din0,
    grp_fu_2529_p_din1,
    grp_fu_2529_p_opcode,
    grp_fu_2529_p_dout0,
    grp_fu_2529_p_ce,
    grp_fu_2533_p_din0,
    grp_fu_2533_p_din1,
    grp_fu_2533_p_dout0,
    grp_fu_2533_p_ce,
    grp_fu_1454_p_din0,
    grp_fu_1454_p_din1,
    grp_fu_1454_p_opcode,
    grp_fu_1454_p_dout0,
    grp_fu_1454_p_ce,
    grp_fu_1462_p_din0,
    grp_fu_1462_p_din1,
    grp_fu_1462_p_dout0,
    grp_fu_1462_p_ce
);

    parameter ap_ST_fsm_pp0_stage0 = 8'd1;
    parameter ap_ST_fsm_pp0_stage1 = 8'd2;
    parameter ap_ST_fsm_pp0_stage2 = 8'd4;
    parameter ap_ST_fsm_pp0_stage3 = 8'd8;
    parameter ap_ST_fsm_pp0_stage4 = 8'd16;
    parameter ap_ST_fsm_pp0_stage5 = 8'd32;
    parameter ap_ST_fsm_pp0_stage6 = 8'd64;
    parameter ap_ST_fsm_pp0_stage7 = 8'd128;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [63:0] minDist;
    input [34:0] sub_ln296;
    output [12:0] rrtVertices_address0;
    output rrtVertices_ce0;
    input [63:0] rrtVertices_q0;
    output [2:0] qRand_address0;
    output qRand_ce0;
    input [63:0] qRand_q0;
    output [11:0] bestIdx_3_out;
    output bestIdx_3_out_ap_vld;
    output [63:0] grp_fu_2529_p_din0;
    output [63:0] grp_fu_2529_p_din1;
    output [1:0] grp_fu_2529_p_opcode;
    input [63:0] grp_fu_2529_p_dout0;
    output grp_fu_2529_p_ce;
    output [63:0] grp_fu_2533_p_din0;
    output [63:0] grp_fu_2533_p_din1;
    input [63:0] grp_fu_2533_p_dout0;
    output grp_fu_2533_p_ce;
    output [63:0] grp_fu_1454_p_din0;
    output [63:0] grp_fu_1454_p_din1;
    output [4:0] grp_fu_1454_p_opcode;
    input [0:0] grp_fu_1454_p_dout0;
    output grp_fu_1454_p_ce;
    output [63:0] grp_fu_1462_p_din0;
    output [63:0] grp_fu_1462_p_din1;
    input [63:0] grp_fu_1462_p_dout0;
    output grp_fu_1462_p_ce;

    reg ap_idle;
    reg rrtVertices_ce0;
    reg qRand_ce0;
    reg bestIdx_3_out_ap_vld;

    (* fsm_encoding = "none" *) reg   [7:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_enable_reg_pp0_iter4;
    reg    ap_enable_reg_pp0_iter5;
    reg    ap_enable_reg_pp0_iter6;
    reg    ap_enable_reg_pp0_iter7;
    reg    ap_enable_reg_pp0_iter8;
    reg    ap_enable_reg_pp0_iter9;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_subdone;
    reg   [0:0] icmp_ln96_reg_497;
    reg    ap_condition_exit_pp0_iter0_stage7;
    wire    ap_loop_exit_ready;
    reg    ap_ready_int;
    wire    ap_block_pp0_stage0_11001;
    reg   [11:0] idx_4_reg_487;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    reg   [11:0] idx_4_reg_487_pp0_iter1_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter2_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter3_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter4_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter5_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter6_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter7_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter8_reg;
    reg   [11:0] idx_4_reg_487_pp0_iter9_reg;
    reg   [34:0] indvar_flatten_load_reg_492;
    wire   [0:0] icmp_ln96_fu_190_p2;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter1_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter2_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter3_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter4_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter5_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter6_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter7_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter8_reg;
    reg   [0:0] icmp_ln96_reg_497_pp0_iter9_reg;
    wire   [0:0] icmp_ln293_fu_204_p2;
    reg   [0:0] icmp_ln293_reg_501;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter1_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter2_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter3_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter4_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter5_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter6_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter7_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter8_reg;
    reg   [0:0] icmp_ln293_reg_501_pp0_iter9_reg;
    wire   [2:0] select_ln96_1_fu_210_p3;
    reg   [2:0] select_ln96_1_reg_508;
    wire   [11:0] select_ln96_3_fu_218_p3;
    reg   [11:0] select_ln96_3_reg_514;
    wire   [9:0] trunc_ln294_fu_226_p1;
    reg   [9:0] trunc_ln294_reg_519;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    reg   [63:0] qRand_load_reg_534;
    reg   [63:0] rrtVertices_load_reg_539;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    reg   [63:0] sub_i9_i_reg_544;
    wire   [63:0] select_ln96_2_fu_298_p3;
    reg   [63:0] select_ln96_2_reg_555;
    reg   [63:0] mul_i10_i_reg_560;
    reg   [63:0] dist_3_reg_565;
    reg   [63:0] d_reg_570;
    reg   [63:0] minDist_7_reg_577;
    reg   [31:0] bestIdx_4_reg_585;
    wire   [0:0] and_ln98_1_fu_395_p2;
    reg   [0:0] and_ln98_1_reg_590;
    wire   [31:0] bestIdx_6_fu_401_p3;
    reg   [31:0] bestIdx_6_reg_595;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage3_subdone;
    reg    ap_condition_exit_pp0_iter9_stage3;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_subdone;
    wire   [63:0] zext_ln293_fu_230_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln294_2_fu_269_p1;
    wire    ap_block_pp0_stage2;
    reg   [63:0] dist_2_fu_68;
    reg   [63:0] ap_sig_allocacmp_dist;
    wire    ap_loop_init;
    reg   [2:0] i_fu_72;
    wire   [2:0] add_ln293_fu_279_p2;
    reg   [31:0] bestIdx_fu_76;
    wire   [31:0] select_ln96_fu_425_p3;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_block_pp0_stage3;
    reg   [63:0] minDist_1_fu_80;
    wire   [63:0] select_ln96_4_fu_419_p3;
    reg   [11:0] idx_fu_84;
    reg   [34:0] indvar_flatten_fu_88;
    wire   [34:0] add_ln96_2_fu_274_p2;
    wire    ap_block_pp0_stage3_01001;
    wire    ap_block_pp0_stage0;
    reg   [63:0] grp_fu_137_p0;
    reg   [63:0] grp_fu_137_p1;
    wire    ap_block_pp0_stage4;
    wire   [11:0] add_ln96_fu_198_p2;
    wire   [12:0] tmp_28_fu_240_p3;
    wire   [12:0] tmp_29_fu_247_p3;
    wire   [12:0] sub_ln294_fu_254_p2;
    wire   [12:0] zext_ln294_fu_260_p1;
    wire   [12:0] add_ln294_fu_263_p2;
    wire   [63:0] bitcast_ln98_fu_319_p1;
    wire   [63:0] bitcast_ln98_1_fu_336_p1;
    wire   [10:0] tmp_361_dup_fu_322_p4;
    wire   [51:0] trunc_ln98_fu_332_p1;
    wire   [0:0] icmp_ln98_1_fu_359_p2;
    wire   [0:0] icmp_ln98_fu_353_p2;
    wire   [10:0] tmp_362_dup_fu_339_p4;
    wire   [51:0] trunc_ln98_2_fu_349_p1;
    wire   [0:0] icmp_ln98_3_fu_377_p2;
    wire   [0:0] icmp_ln98_2_fu_371_p2;
    wire   [0:0] or_ln98_fu_365_p2;
    wire   [0:0] or_ln98_1_fu_383_p2;
    wire   [0:0] and_ln98_fu_389_p2;
    wire   [31:0] zext_ln96_fu_316_p1;
    wire   [63:0] minDist_11_fu_414_p3;
    reg   [1:0] grp_fu_137_opcode;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage4_00001;
    reg    ap_done_reg;
    wire    ap_continue_int;
    reg    ap_done_int;
    reg    ap_loop_exit_ready_pp0_iter1_reg;
    wire    ap_block_pp0_stage7_11001;
    reg    ap_idle_pp0_0to8;
    reg    ap_loop_exit_ready_pp0_iter2_reg;
    reg    ap_loop_exit_ready_pp0_iter3_reg;
    reg    ap_loop_exit_ready_pp0_iter4_reg;
    reg    ap_loop_exit_ready_pp0_iter5_reg;
    reg    ap_loop_exit_ready_pp0_iter6_reg;
    reg    ap_loop_exit_ready_pp0_iter7_reg;
    reg    ap_loop_exit_ready_pp0_iter8_reg;
    reg    ap_loop_exit_ready_pp0_iter9_reg;
    reg   [7:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to9;
    reg    ap_done_pending_pp0;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_enable_pp0;
    wire    ap_start_int;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 8'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter4 = 1'b0;
        #0 ap_enable_reg_pp0_iter5 = 1'b0;
        #0 ap_enable_reg_pp0_iter6 = 1'b0;
        #0 ap_enable_reg_pp0_iter7 = 1'b0;
        #0 ap_enable_reg_pp0_iter8 = 1'b0;
        #0 ap_enable_reg_pp0_iter9 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
        #0 dist_2_fu_68 = 64'd0;
        #0 i_fu_72 = 3'd0;
        #0 bestIdx_fu_76 = 32'd0;
        #0 minDist_1_fu_80 = 64'd0;
        #0 idx_fu_84 = 12'd0;
        #0 indvar_flatten_fu_88 = 35'd0;
        #0 ap_done_reg = 1'b0;
    end

    main_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(ap_start),
        .ap_ready(ap_ready),
        .ap_done(ap_done),
        .ap_start_int(ap_start_int),
        .ap_loop_init(ap_loop_init),
        .ap_ready_int(ap_ready_int),
        .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage7),
        .ap_loop_exit_done(ap_done_int),
        .ap_continue_int(ap_continue_int),
        .ap_done_int(ap_done_int)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_done_reg <= 1'b0;
        end else begin
            if ((ap_continue_int == 1'b1)) begin
                ap_done_reg <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                ap_done_reg <= 1'b1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start_int;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter8 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter9 <= 1'b0;
        end else begin
            if (((1'b1 == ap_condition_exit_pp0_iter9_stage3) | ((1'b0 == ap_block_pp0_stage4_subdone) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
                ap_enable_reg_pp0_iter9 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage7_subdone) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
                ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready_pp0_iter1_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        end
    end

    always @(posedge ap_clk) begin
        if ((((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3)) | ((1'b0 == ap_block_pp0_stage4_subdone) & (ap_loop_exit_ready_pp0_iter8_reg == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage4)))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage7_11001) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            bestIdx_fu_76 <= 32'd0;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln96_reg_497_pp0_iter9_reg == 1'd0))) begin
            bestIdx_fu_76 <= select_ln96_fu_425_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            dist_2_fu_68 <= 64'd0;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_reg_497_pp0_iter2_reg == 1'd0))) begin
            dist_2_fu_68 <= dist_3_reg_565;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                i_fu_72 <= 3'd0;
            end else if (((icmp_ln96_reg_497 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                i_fu_72 <= add_ln293_fu_279_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            idx_fu_84 <= 12'd1;
        end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_fu_190_p2 == 1'd0))) begin
            idx_fu_84 <= select_ln96_3_fu_218_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            if ((ap_loop_init == 1'b1)) begin
                indvar_flatten_fu_88 <= 35'd0;
            end else if (((icmp_ln96_reg_497 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
                indvar_flatten_fu_88 <= add_ln96_2_fu_274_p2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            minDist_1_fu_80 <= minDist;
        end else if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4) & (icmp_ln96_reg_497_pp0_iter9_reg == 1'd0))) begin
            minDist_1_fu_80 <= select_ln96_4_fu_419_p3;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            and_ln98_1_reg_590 <= and_ln98_1_fu_395_p2;
            bestIdx_4_reg_585 <= bestIdx_fu_76;
            bestIdx_6_reg_595 <= bestIdx_6_fu_401_p3;
            rrtVertices_load_reg_539 <= rrtVertices_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            d_reg_570 <= grp_fu_1462_p_dout0;
            icmp_ln293_reg_501 <= icmp_ln293_fu_204_p2;
            icmp_ln293_reg_501_pp0_iter1_reg <= icmp_ln293_reg_501;
            icmp_ln293_reg_501_pp0_iter2_reg <= icmp_ln293_reg_501_pp0_iter1_reg;
            icmp_ln293_reg_501_pp0_iter3_reg <= icmp_ln293_reg_501_pp0_iter2_reg;
            icmp_ln293_reg_501_pp0_iter4_reg <= icmp_ln293_reg_501_pp0_iter3_reg;
            icmp_ln293_reg_501_pp0_iter5_reg <= icmp_ln293_reg_501_pp0_iter4_reg;
            icmp_ln293_reg_501_pp0_iter6_reg <= icmp_ln293_reg_501_pp0_iter5_reg;
            icmp_ln293_reg_501_pp0_iter7_reg <= icmp_ln293_reg_501_pp0_iter6_reg;
            icmp_ln293_reg_501_pp0_iter8_reg <= icmp_ln293_reg_501_pp0_iter7_reg;
            icmp_ln293_reg_501_pp0_iter9_reg <= icmp_ln293_reg_501_pp0_iter8_reg;
            icmp_ln96_reg_497 <= icmp_ln96_fu_190_p2;
            icmp_ln96_reg_497_pp0_iter1_reg <= icmp_ln96_reg_497;
            icmp_ln96_reg_497_pp0_iter2_reg <= icmp_ln96_reg_497_pp0_iter1_reg;
            icmp_ln96_reg_497_pp0_iter3_reg <= icmp_ln96_reg_497_pp0_iter2_reg;
            icmp_ln96_reg_497_pp0_iter4_reg <= icmp_ln96_reg_497_pp0_iter3_reg;
            icmp_ln96_reg_497_pp0_iter5_reg <= icmp_ln96_reg_497_pp0_iter4_reg;
            icmp_ln96_reg_497_pp0_iter6_reg <= icmp_ln96_reg_497_pp0_iter5_reg;
            icmp_ln96_reg_497_pp0_iter7_reg <= icmp_ln96_reg_497_pp0_iter6_reg;
            icmp_ln96_reg_497_pp0_iter8_reg <= icmp_ln96_reg_497_pp0_iter7_reg;
            icmp_ln96_reg_497_pp0_iter9_reg <= icmp_ln96_reg_497_pp0_iter8_reg;
            idx_4_reg_487 <= idx_fu_84;
            idx_4_reg_487_pp0_iter1_reg <= idx_4_reg_487;
            idx_4_reg_487_pp0_iter2_reg <= idx_4_reg_487_pp0_iter1_reg;
            idx_4_reg_487_pp0_iter3_reg <= idx_4_reg_487_pp0_iter2_reg;
            idx_4_reg_487_pp0_iter4_reg <= idx_4_reg_487_pp0_iter3_reg;
            idx_4_reg_487_pp0_iter5_reg <= idx_4_reg_487_pp0_iter4_reg;
            idx_4_reg_487_pp0_iter6_reg <= idx_4_reg_487_pp0_iter5_reg;
            idx_4_reg_487_pp0_iter7_reg <= idx_4_reg_487_pp0_iter6_reg;
            idx_4_reg_487_pp0_iter8_reg <= idx_4_reg_487_pp0_iter7_reg;
            idx_4_reg_487_pp0_iter9_reg <= idx_4_reg_487_pp0_iter8_reg;
            indvar_flatten_load_reg_492 <= indvar_flatten_fu_88;
            mul_i10_i_reg_560 <= grp_fu_2533_p_dout0;
            select_ln96_1_reg_508 <= select_ln96_1_fu_210_p3;
            select_ln96_2_reg_555 <= select_ln96_2_fu_298_p3;
            select_ln96_3_reg_514 <= select_ln96_3_fu_218_p3;
            trunc_ln294_reg_519 <= trunc_ln294_fu_226_p1;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            dist_3_reg_565 <= grp_fu_2529_p_dout0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            minDist_7_reg_577  <= minDist_1_fu_80;
            qRand_load_reg_534 <= qRand_q0;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            sub_i9_i_reg_544 <= grp_fu_2529_p_dout0;
        end
    end

    always @(*) begin
        if (((icmp_ln96_reg_497 == 1'd1) & (1'b0 == ap_block_pp0_stage7_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_condition_exit_pp0_iter0_stage7 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter0_stage7 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_enable_reg_pp0_iter9 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3) & (icmp_ln96_reg_497_pp0_iter9_reg == 1'd1))) begin
            ap_condition_exit_pp0_iter9_stage3 = 1'b1;
        end else begin
            ap_condition_exit_pp0_iter9_stage3 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_done_int = 1'b1;
        end else begin
            ap_done_int = ap_done_reg;
        end
    end

    always @(*) begin
        if (~((ap_loop_exit_ready == 1'b0) & (ap_loop_exit_ready_pp0_iter9_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter8_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter7_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter6_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter5_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter4_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0) & (ap_loop_exit_ready_pp0_iter1_reg == 1'b0))) begin
            ap_done_pending_pp0 = 1'b1;
        end else begin
            ap_done_pending_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start_int;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to8 = 1'b1;
        end else begin
            ap_idle_pp0_0to8 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to9 = 1'b1;
        end else begin
            ap_idle_pp0_1to9 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage7_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            ap_ready_int = 1'b1;
        end else begin
            ap_ready_int = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln96_reg_497_pp0_iter2_reg == 1'd0))) begin
            ap_sig_allocacmp_dist = dist_3_reg_565;
        end else begin
            ap_sig_allocacmp_dist = dist_2_fu_68;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (icmp_ln96_reg_497_pp0_iter9_reg == 1'd1))) begin
            bestIdx_3_out_ap_vld = 1'b1;
        end else begin
            bestIdx_3_out_ap_vld = 1'b0;
        end
    end

    always @(*) begin
        if (((icmp_ln96_reg_497 == 1'd0) & (1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_137_opcode = 2'd1;
        end else if (((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (icmp_ln96_reg_497_pp0_iter2_reg == 1'd0))) begin
            grp_fu_137_opcode = 2'd0;
        end else begin
            grp_fu_137_opcode = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_137_p0 = select_ln96_2_reg_555;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_137_p0 = rrtVertices_load_reg_539;
        end else begin
            grp_fu_137_p0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_137_p1 = mul_i10_i_reg_560;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_137_p1 = qRand_load_reg_534;
        end else begin
            grp_fu_137_p1 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            qRand_ce0 = 1'b1;
        end else begin
            qRand_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            rrtVertices_ce0 = 1'b1;
        end else begin
            rrtVertices_ce0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start_int == 1'b0) & (ap_done_pending_pp0 == 1'b0) & (ap_idle_pp0_1to9 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if (((ap_idle_pp0_0to8 == 1'b1) & (1'b1 == ap_condition_exit_pp0_iter9_stage3))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln293_fu_279_p2 = (select_ln96_1_reg_508 + 3'd1);

    assign add_ln294_fu_263_p2 = (sub_ln294_fu_254_p2 + zext_ln294_fu_260_p1);

    assign add_ln96_2_fu_274_p2 = (indvar_flatten_load_reg_492 + 35'd1);

    assign add_ln96_fu_198_p2 = (idx_fu_84 + 12'd1);

    assign and_ln98_1_fu_395_p2 = (grp_fu_1454_p_dout0 & and_ln98_fu_389_p2);

    assign and_ln98_fu_389_p2 = (or_ln98_fu_365_p2 & or_ln98_1_fu_383_p2);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_01001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage7;

    assign bestIdx_3_out = bestIdx_6_fu_401_p3[11:0];

    assign bestIdx_6_fu_401_p3 = ((and_ln98_1_fu_395_p2[0:0] == 1'b1) ? zext_ln96_fu_316_p1 : bestIdx_fu_76);

    assign bitcast_ln98_1_fu_336_p1 = minDist_7_reg_577;

    assign bitcast_ln98_fu_319_p1 = d_reg_570;

    assign grp_fu_1454_p_ce = 1'b1;

    assign grp_fu_1454_p_din0 = d_reg_570;

    assign grp_fu_1454_p_din1 = minDist_1_fu_80;

    assign grp_fu_1454_p_opcode = 5'd4;

    assign grp_fu_1462_p_ce = 1'b1;

    assign grp_fu_1462_p_din0 = 64'd0;

    assign grp_fu_1462_p_din1 = ap_sig_allocacmp_dist;

    assign grp_fu_2529_p_ce = 1'b1;

    assign grp_fu_2529_p_din0 = grp_fu_137_p0;

    assign grp_fu_2529_p_din1 = grp_fu_137_p1;

    assign grp_fu_2529_p_opcode = grp_fu_137_opcode;

    assign grp_fu_2533_p_ce = 1'b1;

    assign grp_fu_2533_p_din0 = sub_i9_i_reg_544;

    assign grp_fu_2533_p_din1 = sub_i9_i_reg_544;

    assign icmp_ln293_fu_204_p2 = ((i_fu_72 == 3'd6) ? 1'b1 : 1'b0);

    assign icmp_ln96_fu_190_p2 = ((indvar_flatten_fu_88 == sub_ln296) ? 1'b1 : 1'b0);

    assign icmp_ln98_1_fu_359_p2 = ((trunc_ln98_fu_332_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln98_2_fu_371_p2 = ((tmp_362_dup_fu_339_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign icmp_ln98_3_fu_377_p2 = ((trunc_ln98_2_fu_349_p1 == 52'd0) ? 1'b1 : 1'b0);

    assign icmp_ln98_fu_353_p2 = ((tmp_361_dup_fu_322_p4 != 11'd2047) ? 1'b1 : 1'b0);

    assign minDist_11_fu_414_p3 = ((and_ln98_1_reg_590[0:0] == 1'b1) ? d_reg_570 : minDist_7_reg_577);

    assign or_ln98_1_fu_383_p2 = (icmp_ln98_3_fu_377_p2 | icmp_ln98_2_fu_371_p2);

    assign or_ln98_fu_365_p2 = (icmp_ln98_fu_353_p2 | icmp_ln98_1_fu_359_p2);

    assign qRand_address0 = zext_ln293_fu_230_p1;

    assign rrtVertices_address0 = zext_ln294_2_fu_269_p1;

    assign select_ln96_1_fu_210_p3 = ((icmp_ln293_fu_204_p2[0:0] == 1'b1) ? 3'd0 : i_fu_72);

    assign select_ln96_2_fu_298_p3 = ((icmp_ln293_reg_501_pp0_iter1_reg[0:0] == 1'b1) ? 64'd0 : ap_sig_allocacmp_dist);

    assign select_ln96_3_fu_218_p3 = ((icmp_ln293_fu_204_p2[0:0] == 1'b1) ? add_ln96_fu_198_p2 : idx_fu_84);

    assign select_ln96_4_fu_419_p3 = ((icmp_ln293_reg_501_pp0_iter9_reg[0:0] == 1'b1) ? minDist_11_fu_414_p3 : minDist_7_reg_577);

    assign select_ln96_fu_425_p3 = ((icmp_ln293_reg_501_pp0_iter9_reg[0:0] == 1'b1) ? bestIdx_6_reg_595 : bestIdx_4_reg_585);

    assign sub_ln294_fu_254_p2 = (tmp_28_fu_240_p3 - tmp_29_fu_247_p3);

    assign tmp_28_fu_240_p3 = {{trunc_ln294_reg_519}, {3'd0}};

    assign tmp_29_fu_247_p3 = {{select_ln96_3_reg_514}, {1'd0}};

    assign tmp_361_dup_fu_322_p4 = {{bitcast_ln98_fu_319_p1[62:52]}};

    assign tmp_362_dup_fu_339_p4 = {{bitcast_ln98_1_fu_336_p1[62:52]}};

    assign trunc_ln294_fu_226_p1 = select_ln96_3_fu_218_p3[9:0];

    assign trunc_ln98_2_fu_349_p1 = bitcast_ln98_1_fu_336_p1[51:0];

    assign trunc_ln98_fu_332_p1 = bitcast_ln98_fu_319_p1[51:0];

    assign zext_ln293_fu_230_p1 = select_ln96_1_fu_210_p3;

    assign zext_ln294_2_fu_269_p1 = add_ln294_fu_263_p2;

    assign zext_ln294_fu_260_p1 = select_ln96_1_reg_508;

    assign zext_ln96_fu_316_p1 = idx_4_reg_487_pp0_iter9_reg;

endmodule  //main_planRRT_Pipeline_VITIS_LOOP_96_2_VITIS_LOOP_293_1
