/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_blockDescToBoundingBox_double_s (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    H_offset,
    dim_0_0_val,
    dim_0_1_val,
    dim_0_2_val,
    corners_address0,
    corners_ce0,
    corners_we0,
    corners_d0,
    corners_address1,
    corners_ce1,
    corners_we1,
    corners_d1,
    l_TColl_0_0_0_constprop,
    l_TColl_0_0_1_constprop,
    l_TColl_0_0_2_constprop,
    l_TColl_0_0_3_constprop,
    l_TColl_1_0_0_constprop,
    l_TColl_1_0_1_constprop,
    l_TColl_1_0_2_constprop,
    l_TColl_1_0_3_constprop,
    l_TColl_2_0_0_constprop,
    l_TColl_2_0_1_constprop,
    l_TColl_2_0_2_constprop,
    l_TColl_2_0_3_constprop,
    l_TColl_0_1_0_constprop,
    l_TColl_0_1_1_constprop,
    l_TColl_0_1_2_constprop,
    l_TColl_0_1_3_constprop,
    l_TColl_1_1_0_constprop,
    l_TColl_1_1_1_constprop,
    l_TColl_1_1_2_constprop,
    l_TColl_1_1_3_constprop,
    l_TColl_2_1_0_constprop,
    l_TColl_2_1_1_constprop,
    l_TColl_2_1_2_constprop,
    l_TColl_2_1_3_constprop,
    l_TColl_0_2_0_constprop,
    l_TColl_0_2_1_constprop,
    l_TColl_0_2_2_constprop,
    l_TColl_0_2_3_constprop,
    l_TColl_1_2_0_constprop,
    l_TColl_1_2_1_constprop,
    l_TColl_1_2_2_constprop,
    l_TColl_1_2_3_constprop,
    l_TColl_2_2_0_constprop,
    l_TColl_2_2_1_constprop,
    l_TColl_2_2_2_constprop,
    l_TColl_2_2_3_constprop,
    l_TColl_0_3_0_constprop,
    l_TColl_0_3_1_constprop,
    l_TColl_0_3_2_constprop,
    l_TColl_0_3_3_constprop,
    l_TColl_1_3_0_constprop,
    l_TColl_1_3_1_constprop,
    l_TColl_1_3_2_constprop,
    l_TColl_1_3_3_constprop,
    l_TColl_2_3_0_constprop,
    l_TColl_2_3_1_constprop,
    l_TColl_2_3_2_constprop,
    l_TColl_2_3_3_constprop
);

    parameter ap_ST_fsm_pp0_stage0 = 14'd1;
    parameter ap_ST_fsm_pp0_stage1 = 14'd2;
    parameter ap_ST_fsm_pp0_stage2 = 14'd4;
    parameter ap_ST_fsm_pp0_stage3 = 14'd8;
    parameter ap_ST_fsm_pp0_stage4 = 14'd16;
    parameter ap_ST_fsm_pp0_stage5 = 14'd32;
    parameter ap_ST_fsm_pp0_stage6 = 14'd64;
    parameter ap_ST_fsm_pp0_stage7 = 14'd128;
    parameter ap_ST_fsm_pp0_stage8 = 14'd256;
    parameter ap_ST_fsm_pp0_stage9 = 14'd512;
    parameter ap_ST_fsm_pp0_stage10 = 14'd1024;
    parameter ap_ST_fsm_pp0_stage11 = 14'd2048;
    parameter ap_ST_fsm_pp0_stage12 = 14'd4096;
    parameter ap_ST_fsm_pp0_stage13 = 14'd8192;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    input [1:0] H_offset;
    input [63:0] dim_0_0_val;
    input [63:0] dim_0_1_val;
    input [63:0] dim_0_2_val;
    output [6:0] corners_address0;
    output corners_ce0;
    output corners_we0;
    output [63:0] corners_d0;
    output [6:0] corners_address1;
    output corners_ce1;
    output corners_we1;
    output [63:0] corners_d1;
    input [63:0] l_TColl_0_0_0_constprop;
    input [63:0] l_TColl_0_0_1_constprop;
    input [63:0] l_TColl_0_0_2_constprop;
    input [63:0] l_TColl_0_0_3_constprop;
    input [63:0] l_TColl_1_0_0_constprop;
    input [63:0] l_TColl_1_0_1_constprop;
    input [63:0] l_TColl_1_0_2_constprop;
    input [63:0] l_TColl_1_0_3_constprop;
    input [63:0] l_TColl_2_0_0_constprop;
    input [63:0] l_TColl_2_0_1_constprop;
    input [63:0] l_TColl_2_0_2_constprop;
    input [63:0] l_TColl_2_0_3_constprop;
    input [63:0] l_TColl_0_1_0_constprop;
    input [63:0] l_TColl_0_1_1_constprop;
    input [63:0] l_TColl_0_1_2_constprop;
    input [63:0] l_TColl_0_1_3_constprop;
    input [63:0] l_TColl_1_1_0_constprop;
    input [63:0] l_TColl_1_1_1_constprop;
    input [63:0] l_TColl_1_1_2_constprop;
    input [63:0] l_TColl_1_1_3_constprop;
    input [63:0] l_TColl_2_1_0_constprop;
    input [63:0] l_TColl_2_1_1_constprop;
    input [63:0] l_TColl_2_1_2_constprop;
    input [63:0] l_TColl_2_1_3_constprop;
    input [63:0] l_TColl_0_2_0_constprop;
    input [63:0] l_TColl_0_2_1_constprop;
    input [63:0] l_TColl_0_2_2_constprop;
    input [63:0] l_TColl_0_2_3_constprop;
    input [63:0] l_TColl_1_2_0_constprop;
    input [63:0] l_TColl_1_2_1_constprop;
    input [63:0] l_TColl_1_2_2_constprop;
    input [63:0] l_TColl_1_2_3_constprop;
    input [63:0] l_TColl_2_2_0_constprop;
    input [63:0] l_TColl_2_2_1_constprop;
    input [63:0] l_TColl_2_2_2_constprop;
    input [63:0] l_TColl_2_2_3_constprop;
    input [63:0] l_TColl_0_3_0_constprop;
    input [63:0] l_TColl_0_3_1_constprop;
    input [63:0] l_TColl_0_3_2_constprop;
    input [63:0] l_TColl_0_3_3_constprop;
    input [63:0] l_TColl_1_3_0_constprop;
    input [63:0] l_TColl_1_3_1_constprop;
    input [63:0] l_TColl_1_3_2_constprop;
    input [63:0] l_TColl_1_3_3_constprop;
    input [63:0] l_TColl_2_3_0_constprop;
    input [63:0] l_TColl_2_3_1_constprop;
    input [63:0] l_TColl_2_3_2_constprop;
    input [63:0] l_TColl_2_3_3_constprop;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[6:0] corners_address0;
    reg corners_ce0;
    reg corners_we0;
    reg[63:0] corners_d0;
    reg[6:0] corners_address1;
    reg corners_ce1;
    reg corners_we1;
    reg[63:0] corners_d1;

    (* fsm_encoding = "none" *) reg   [13:0] ap_CS_fsm;
    wire    ap_CS_fsm_pp0_stage0;
    reg    ap_enable_reg_pp0_iter0;
    reg    ap_enable_reg_pp0_iter1;
    reg    ap_enable_reg_pp0_iter2;
    reg    ap_enable_reg_pp0_iter3;
    reg    ap_idle_pp0;
    wire    ap_CS_fsm_pp0_stage13;
    wire    ap_block_pp0_stage13_subdone;
    wire   [63:0] grp_fu_431_p2;
    reg   [63:0] reg_446;
    wire    ap_CS_fsm_pp0_stage7;
    wire    ap_block_pp0_stage7_11001;
    wire    ap_block_pp0_stage0_11001;
    reg   [63:0] reg_453;
    wire    ap_CS_fsm_pp0_stage8;
    wire    ap_block_pp0_stage8_11001;
    wire    ap_CS_fsm_pp0_stage1;
    wire    ap_block_pp0_stage1_11001;
    wire   [63:0] grp_fu_419_p2;
    reg   [63:0] reg_460;
    wire    ap_CS_fsm_pp0_stage4;
    wire    ap_block_pp0_stage4_11001;
    wire    ap_CS_fsm_pp0_stage5;
    wire    ap_block_pp0_stage5_11001;
    wire   [63:0] grp_fu_423_p2;
    reg   [63:0] reg_468;
    wire   [63:0] grp_fu_427_p2;
    reg   [63:0] reg_475;
    reg   [63:0] reg_481;
    wire    ap_CS_fsm_pp0_stage6;
    wire    ap_block_pp0_stage6_11001;
    reg   [63:0] reg_488;
    reg   [63:0] reg_494;
    reg   [63:0] reg_500;
    wire    ap_CS_fsm_pp0_stage10;
    wire    ap_block_pp0_stage10_11001;
    wire    ap_CS_fsm_pp0_stage11;
    wire    ap_block_pp0_stage11_11001;
    reg   [63:0] reg_507;
    reg   [63:0] reg_513;
    wire    ap_CS_fsm_pp0_stage9;
    wire    ap_block_pp0_stage9_11001;
    wire    ap_CS_fsm_pp0_stage12;
    wire    ap_block_pp0_stage12_11001;
    reg   [63:0] reg_519;
    wire    ap_block_pp0_stage13_11001;
    reg   [63:0] reg_524;
    reg   [63:0] reg_529;
    reg   [1:0] H_offset_read_reg_1163;
    wire   [6:0] mul_ln50_fu_538_p2;
    reg   [6:0] mul_ln50_reg_1176;
    reg   [6:0] mul_ln50_reg_1176_pp0_iter1_reg;
    reg   [6:0] mul_ln50_reg_1176_pp0_iter2_reg;
    reg   [6:0] mul_ln50_reg_1176_pp0_iter3_reg;
    wire   [63:0] tmp_fu_565_p6;
    reg   [63:0] tmp_reg_1206;
    wire   [63:0] tmp_s_fu_595_p6;
    reg   [63:0] tmp_s_reg_1211;
    wire   [63:0] tmp_314_fu_625_p6;
    reg   [63:0] tmp_314_reg_1216;
    reg   [63:0] tmp_314_reg_1216_pp0_iter1_reg;
    reg   [63:0] dim_0_0_val_read_reg_1222;
    wire   [63:0] tmp_307_fu_676_p6;
    reg   [63:0] tmp_307_reg_1228;
    wire   [63:0] tmp_308_fu_705_p6;
    reg   [63:0] tmp_308_reg_1233;
    wire   [63:0] tmp_315_fu_734_p6;
    reg   [63:0] tmp_315_reg_1238;
    reg   [63:0] tmp_315_reg_1238_pp0_iter1_reg;
    wire   [63:0] tmp_316_fu_764_p6;
    reg   [63:0] tmp_316_reg_1243;
    reg   [63:0] tmp_316_reg_1243_pp0_iter1_reg;
    reg   [63:0] dim_0_1_val_read_reg_1249;
    wire    ap_CS_fsm_pp0_stage2;
    wire    ap_block_pp0_stage2_11001;
    wire   [63:0] tmp_309_fu_794_p6;
    reg   [63:0] tmp_309_reg_1255;
    wire   [63:0] tmp_310_fu_823_p6;
    reg   [63:0] tmp_310_reg_1260;
    wire   [63:0] tmp_311_fu_852_p6;
    reg   [63:0] tmp_311_reg_1265;
    wire    ap_CS_fsm_pp0_stage3;
    wire    ap_block_pp0_stage3_11001;
    wire   [63:0] tmp_312_fu_881_p6;
    reg   [63:0] tmp_312_reg_1270;
    reg   [63:0] dim_0_2_val_read_reg_1275;
    wire   [63:0] tmp_313_fu_910_p6;
    reg   [63:0] tmp_313_reg_1281;
    wire   [63:0] grp_fu_436_p2;
    reg   [63:0] mul6_reg_1286;
    reg   [63:0] mul4_reg_1291;
    reg   [63:0] mul5_reg_1296;
    reg   [63:0] mul7_reg_1301;
    reg   [63:0] mul8_reg_1306;
    reg   [63:0] mul9_reg_1311;
    reg   [63:0] mul1_reg_1316;
    reg   [63:0] xL_1_reg_1321;
    reg   [63:0] yL_reg_1326;
    reg   [63:0] yL_1_reg_1332;
    reg   [63:0] yL_2_reg_1337;
    reg   [63:0] zL_reg_1343;
    reg   [63:0] zL_reg_1343_pp0_iter2_reg;
    reg   [63:0] zL_1_reg_1348;
    reg   [63:0] zL_1_reg_1348_pp0_iter2_reg;
    reg   [63:0] zL_2_reg_1353;
    reg   [63:0] zL_2_reg_1353_pp0_iter2_reg;
    reg   [63:0] sub3_reg_1358;
    reg   [63:0] add67_2_reg_1363;
    reg   [63:0] sub112_1_reg_1368;
    reg   [63:0] sub112_2_reg_1373;
    reg   [63:0] add5_reg_1378;
    reg   [63:0] add158_1_reg_1383;
    reg   [63:0] add158_2_reg_1388;
    reg   [63:0] sub7_reg_1393;
    reg   [63:0] sub204_1_reg_1398;
    reg   [63:0] sub204_2_reg_1403;
    reg   [63:0] sub138_1_reg_1408;
    reg   [63:0] add6_reg_1413;
    reg   [63:0] add161_2_reg_1418;
    reg    ap_enable_reg_pp0_iter0_reg;
    wire    ap_block_pp0_stage9_subdone;
    reg   [63:0] ap_port_reg_dim_0_0_val;
    reg   [63:0] ap_port_reg_dim_0_1_val;
    reg   [63:0] ap_port_reg_dim_0_2_val;
    wire   [63:0] zext_ln50_1_fu_544_p1;
    wire    ap_block_pp0_stage0;
    wire   [63:0] zext_ln50_2_fu_645_p1;
    wire    ap_block_pp0_stage1;
    wire   [63:0] zext_ln50_3_fu_655_p1;
    wire   [63:0] zext_ln51_fu_928_p1;
    wire    ap_block_pp0_stage10;
    wire   [63:0] zext_ln51_1_fu_938_p1;
    wire   [63:0] zext_ln51_2_fu_948_p1;
    wire    ap_block_pp0_stage11;
    wire   [63:0] zext_ln52_fu_958_p1;
    wire   [63:0] zext_ln52_1_fu_968_p1;
    wire    ap_block_pp0_stage12;
    wire   [63:0] zext_ln52_2_fu_978_p1;
    wire   [63:0] zext_ln53_fu_988_p1;
    wire    ap_block_pp0_stage13;
    wire   [63:0] zext_ln53_1_fu_998_p1;
    wire   [63:0] zext_ln53_2_fu_1008_p1;
    wire   [63:0] zext_ln54_fu_1018_p1;
    wire    ap_block_pp0_stage2;
    wire   [63:0] zext_ln54_1_fu_1028_p1;
    wire   [63:0] zext_ln54_2_fu_1038_p1;
    wire    ap_block_pp0_stage3;
    wire   [63:0] zext_ln55_fu_1048_p1;
    wire   [63:0] zext_ln55_1_fu_1058_p1;
    wire    ap_block_pp0_stage4;
    wire   [63:0] zext_ln55_2_fu_1068_p1;
    wire   [63:0] zext_ln56_fu_1078_p1;
    wire    ap_block_pp0_stage5;
    wire   [63:0] zext_ln56_1_fu_1088_p1;
    wire   [63:0] zext_ln56_2_fu_1098_p1;
    wire    ap_block_pp0_stage6;
    wire   [63:0] zext_ln57_fu_1108_p1;
    wire   [63:0] zext_ln57_1_fu_1118_p1;
    wire    ap_block_pp0_stage7;
    wire   [63:0] zext_ln57_2_fu_1128_p1;
    wire   [63:0] zext_ln58_fu_1138_p1;
    wire    ap_block_pp0_stage8;
    wire   [63:0] zext_ln58_1_fu_1148_p1;
    wire   [63:0] zext_ln58_2_fu_1158_p1;
    wire    ap_block_pp0_stage9;
    reg   [63:0] grp_fu_419_p0;
    reg   [63:0] grp_fu_419_p1;
    reg   [63:0] grp_fu_423_p0;
    reg   [63:0] grp_fu_423_p1;
    reg   [63:0] grp_fu_427_p0;
    reg   [63:0] grp_fu_427_p1;
    reg   [63:0] grp_fu_431_p0;
    reg   [63:0] grp_fu_431_p1;
    reg   [63:0] grp_fu_436_p0;
    reg   [63:0] grp_fu_436_p1;
    wire   [1:0] mul_ln50_fu_538_p0;
    wire   [5:0] mul_ln50_fu_538_p1;
    wire   [6:0] add_ln50_fu_640_p2;
    wire   [6:0] add_ln50_1_fu_650_p2;
    wire   [6:0] add_ln51_fu_923_p2;
    wire   [6:0] add_ln51_1_fu_933_p2;
    wire   [6:0] add_ln51_2_fu_943_p2;
    wire   [6:0] add_ln52_fu_953_p2;
    wire   [6:0] add_ln52_1_fu_963_p2;
    wire   [6:0] add_ln52_2_fu_973_p2;
    wire   [6:0] add_ln53_fu_983_p2;
    wire   [6:0] add_ln53_1_fu_993_p2;
    wire   [6:0] add_ln53_2_fu_1003_p2;
    wire   [6:0] add_ln54_fu_1013_p2;
    wire   [6:0] add_ln54_1_fu_1023_p2;
    wire   [6:0] add_ln54_2_fu_1033_p2;
    wire   [6:0] add_ln55_fu_1043_p2;
    wire   [6:0] add_ln55_1_fu_1053_p2;
    wire   [6:0] add_ln55_2_fu_1063_p2;
    wire   [6:0] add_ln56_fu_1073_p2;
    wire   [6:0] add_ln56_1_fu_1083_p2;
    wire   [6:0] add_ln56_2_fu_1093_p2;
    wire   [6:0] add_ln57_fu_1103_p2;
    wire   [6:0] add_ln57_1_fu_1113_p2;
    wire   [6:0] add_ln57_2_fu_1123_p2;
    wire   [6:0] add_ln58_fu_1133_p2;
    wire   [6:0] add_ln58_1_fu_1143_p2;
    wire   [6:0] add_ln58_2_fu_1153_p2;
    reg   [1:0] grp_fu_419_opcode;
    wire    ap_block_pp0_stage1_00001;
    wire    ap_block_pp0_stage2_00001;
    wire    ap_block_pp0_stage8_00001;
    wire    ap_block_pp0_stage9_00001;
    wire    ap_block_pp0_stage10_00001;
    wire    ap_block_pp0_stage3_00001;
    wire    ap_block_pp0_stage5_00001;
    wire    ap_block_pp0_stage7_00001;
    wire    ap_block_pp0_stage13_00001;
    wire    ap_block_pp0_stage11_00001;
    wire    ap_block_pp0_stage4_00001;
    wire    ap_block_pp0_stage6_00001;
    wire    ap_block_pp0_stage12_00001;
    wire    ap_block_pp0_stage0_00001;
    reg   [1:0] grp_fu_423_opcode;
    reg   [1:0] grp_fu_427_opcode;
    reg   [13:0] ap_NS_fsm;
    wire    ap_block_pp0_stage0_subdone;
    reg    ap_idle_pp0_1to3;
    wire    ap_block_pp0_stage1_subdone;
    wire    ap_block_pp0_stage2_subdone;
    wire    ap_block_pp0_stage3_subdone;
    wire    ap_block_pp0_stage4_subdone;
    wire    ap_block_pp0_stage5_subdone;
    wire    ap_block_pp0_stage6_subdone;
    wire    ap_block_pp0_stage7_subdone;
    wire    ap_block_pp0_stage8_subdone;
    reg    ap_idle_pp0_0to2;
    reg    ap_reset_idle_pp0;
    wire    ap_block_pp0_stage10_subdone;
    wire    ap_block_pp0_stage11_subdone;
    wire    ap_block_pp0_stage12_subdone;
    wire    ap_enable_pp0;
    wire   [6:0] mul_ln50_fu_538_p00;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 14'd1;
        #0 ap_enable_reg_pp0_iter1 = 1'b0;
        #0 ap_enable_reg_pp0_iter2 = 1'b0;
        #0 ap_enable_reg_pp0_iter3 = 1'b0;
        #0 ap_enable_reg_pp0_iter0_reg = 1'b0;
    end

    main_dadddsub_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_x_U873 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_419_p0),
        .din1(grp_fu_419_p1),
        .opcode(grp_fu_419_opcode),
        .ce(1'b1),
        .dout(grp_fu_419_p2)
    );

    main_dadddsub_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_x_U874 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_423_p0),
        .din1(grp_fu_423_p1),
        .opcode(grp_fu_423_opcode),
        .ce(1'b1),
        .dout(grp_fu_423_p2)
    );

    main_dadddsub_64ns_64ns_64_7_full_dsp_1_x #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dadddsub_64ns_64ns_64_7_full_dsp_1_x_U875 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_427_p0),
        .din1(grp_fu_427_p1),
        .opcode(grp_fu_427_opcode),
        .ce(1'b1),
        .dout(grp_fu_427_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U876 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_431_p0),
        .din1(grp_fu_431_p1),
        .ce(1'b1),
        .dout(grp_fu_431_p2)
    );

    main_dmul_64ns_64ns_64_7_max_dsp_1 #(
        .ID(1),
        .NUM_STAGE(7),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .dout_WIDTH(64)
    ) dmul_64ns_64ns_64_7_max_dsp_1_U877 (
        .clk(ap_clk),
        .reset(ap_rst),
        .din0(grp_fu_436_p0),
        .din1(grp_fu_436_p1),
        .ce(1'b1),
        .dout(grp_fu_436_p2)
    );

    main_mul_2ns_6ns_7_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(2),
        .din1_WIDTH(6),
        .dout_WIDTH(7)
    ) mul_2ns_6ns_7_1_1_U878 (
        .din0(mul_ln50_fu_538_p0),
        .din1(mul_ln50_fu_538_p1),
        .dout(mul_ln50_fu_538_p2)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U879 (
        .din0(l_TColl_0_0_0_constprop),
        .din1(l_TColl_0_0_1_constprop),
        .din2(l_TColl_0_0_2_constprop),
        .din3(l_TColl_0_0_3_constprop),
        .din4(H_offset),
        .dout(tmp_fu_565_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U880 (
        .din0(l_TColl_1_0_0_constprop),
        .din1(l_TColl_1_0_1_constprop),
        .din2(l_TColl_1_0_2_constprop),
        .din3(l_TColl_1_0_3_constprop),
        .din4(H_offset),
        .dout(tmp_s_fu_595_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U881 (
        .din0(l_TColl_0_3_0_constprop),
        .din1(l_TColl_0_3_1_constprop),
        .din2(l_TColl_0_3_2_constprop),
        .din3(l_TColl_0_3_3_constprop),
        .din4(H_offset),
        .dout(tmp_314_fu_625_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U882 (
        .din0(l_TColl_2_0_0_constprop),
        .din1(l_TColl_2_0_1_constprop),
        .din2(l_TColl_2_0_2_constprop),
        .din3(l_TColl_2_0_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_307_fu_676_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U883 (
        .din0(l_TColl_0_1_0_constprop),
        .din1(l_TColl_0_1_1_constprop),
        .din2(l_TColl_0_1_2_constprop),
        .din3(l_TColl_0_1_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_308_fu_705_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U884 (
        .din0(l_TColl_1_3_0_constprop),
        .din1(l_TColl_1_3_1_constprop),
        .din2(l_TColl_1_3_2_constprop),
        .din3(l_TColl_1_3_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_315_fu_734_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U885 (
        .din0(l_TColl_2_3_0_constprop),
        .din1(l_TColl_2_3_1_constprop),
        .din2(l_TColl_2_3_2_constprop),
        .din3(l_TColl_2_3_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_316_fu_764_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U886 (
        .din0(l_TColl_1_1_0_constprop),
        .din1(l_TColl_1_1_1_constprop),
        .din2(l_TColl_1_1_2_constprop),
        .din3(l_TColl_1_1_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_309_fu_794_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U887 (
        .din0(l_TColl_2_1_0_constprop),
        .din1(l_TColl_2_1_1_constprop),
        .din2(l_TColl_2_1_2_constprop),
        .din3(l_TColl_2_1_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_310_fu_823_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U888 (
        .din0(l_TColl_0_2_0_constprop),
        .din1(l_TColl_0_2_1_constprop),
        .din2(l_TColl_0_2_2_constprop),
        .din3(l_TColl_0_2_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_311_fu_852_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U889 (
        .din0(l_TColl_1_2_0_constprop),
        .din1(l_TColl_1_2_1_constprop),
        .din2(l_TColl_1_2_2_constprop),
        .din3(l_TColl_1_2_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_312_fu_881_p6)
    );

    main_mux_4_2_64_1_1 #(
        .ID(1),
        .NUM_STAGE(1),
        .din0_WIDTH(64),
        .din1_WIDTH(64),
        .din2_WIDTH(64),
        .din3_WIDTH(64),
        .din4_WIDTH(2),
        .dout_WIDTH(64)
    ) mux_4_2_64_1_1_U890 (
        .din0(l_TColl_2_2_0_constprop),
        .din1(l_TColl_2_2_1_constprop),
        .din2(l_TColl_2_2_2_constprop),
        .din3(l_TColl_2_2_3_constprop),
        .din4(H_offset_read_reg_1163),
        .dout(tmp_313_fu_910_p6)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter0_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
                ap_enable_reg_pp0_iter0_reg <= ap_start;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end else begin
            if (((1'b0 == ap_block_pp0_stage9_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                ap_enable_reg_pp0_iter3 <= 1'b0;
            end else if (((1'b0 == ap_block_pp0_stage13_subdone) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
                ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            H_offset_read_reg_1163 <= H_offset;
            mul_ln50_reg_1176 <= mul_ln50_fu_538_p2;
            mul_ln50_reg_1176_pp0_iter1_reg <= mul_ln50_reg_1176;
            mul_ln50_reg_1176_pp0_iter2_reg <= mul_ln50_reg_1176_pp0_iter1_reg;
            mul_ln50_reg_1176_pp0_iter3_reg <= mul_ln50_reg_1176_pp0_iter2_reg;
            tmp_314_reg_1216 <= tmp_314_fu_625_p6;
            tmp_314_reg_1216_pp0_iter1_reg <= tmp_314_reg_1216;
            tmp_reg_1206 <= tmp_fu_565_p6;
            tmp_s_reg_1211 <= tmp_s_fu_595_p6;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            add158_1_reg_1383 <= grp_fu_423_p2;
            add158_2_reg_1388 <= grp_fu_427_p2;
            add5_reg_1378 <= grp_fu_419_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            add161_2_reg_1418 <= grp_fu_427_p2;
            add6_reg_1413 <= grp_fu_419_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            add67_2_reg_1363  <= grp_fu_419_p2;
            sub112_1_reg_1368 <= grp_fu_423_p2;
            sub112_2_reg_1373 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_port_reg_dim_0_0_val <= dim_0_0_val;
            ap_port_reg_dim_0_1_val <= dim_0_1_val;
            ap_port_reg_dim_0_2_val <= dim_0_2_val;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            dim_0_0_val_read_reg_1222 <= ap_port_reg_dim_0_0_val;
            tmp_307_reg_1228 <= tmp_307_fu_676_p6;
            tmp_308_reg_1233 <= tmp_308_fu_705_p6;
            tmp_315_reg_1238 <= tmp_315_fu_734_p6;
            tmp_315_reg_1238_pp0_iter1_reg <= tmp_315_reg_1238;
            tmp_316_reg_1243 <= tmp_316_fu_764_p6;
            tmp_316_reg_1243_pp0_iter1_reg <= tmp_316_reg_1243;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            dim_0_1_val_read_reg_1249 <= ap_port_reg_dim_0_1_val;
            tmp_309_reg_1255 <= tmp_309_fu_794_p6;
            tmp_310_reg_1260 <= tmp_310_fu_823_p6;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            dim_0_2_val_read_reg_1275 <= ap_port_reg_dim_0_2_val;
            tmp_313_reg_1281 <= tmp_313_fu_910_p6;
            zL_2_reg_1353_pp0_iter2_reg <= zL_2_reg_1353;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            mul1_reg_1316 <= grp_fu_431_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            mul4_reg_1291 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            mul5_reg_1296 <= grp_fu_431_p2;
            mul7_reg_1301 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            mul6_reg_1286 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            mul8_reg_1306 <= grp_fu_431_p2;
            mul9_reg_1311 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_446 <= grp_fu_431_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_453 <= grp_fu_431_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_460 <= grp_fu_419_p2;
            reg_468 <= grp_fu_423_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            reg_475 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_481 <= grp_fu_419_p2;
            reg_488 <= grp_fu_423_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            reg_494 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            reg_500 <= grp_fu_419_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            reg_507 <= grp_fu_423_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)))) begin
            reg_513 <= grp_fu_419_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            reg_519 <= grp_fu_423_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)))) begin
            reg_524 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if ((((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            reg_529 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            sub138_1_reg_1408 <= grp_fu_423_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            sub204_1_reg_1398 <= grp_fu_423_p2;
            sub204_2_reg_1403 <= grp_fu_427_p2;
            sub7_reg_1393 <= grp_fu_419_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            sub3_reg_1358 <= grp_fu_427_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            tmp_311_reg_1265 <= tmp_311_fu_852_p6;
            tmp_312_reg_1270 <= tmp_312_fu_881_p6;
            zL_1_reg_1348_pp0_iter2_reg <= zL_1_reg_1348;
            zL_reg_1343_pp0_iter2_reg <= zL_reg_1343;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            xL_1_reg_1321 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            yL_1_reg_1332 <= grp_fu_431_p2;
            yL_2_reg_1337 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            yL_reg_1326 <= grp_fu_436_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            zL_1_reg_1348 <= grp_fu_436_p2;
            zL_reg_1343   <= grp_fu_431_p2;
        end
    end

    always @(posedge ap_clk) begin
        if (((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            zL_2_reg_1353 <= grp_fu_431_p2;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0 = ap_start;
        end else begin
            ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
        end
    end

    always @(*) begin
        if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start == 1'b0))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0 = 1'b1;
        end else begin
            ap_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
            ap_idle_pp0_0to2 = 1'b1;
        end else begin
            ap_idle_pp0_0to2 = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
            ap_idle_pp0_1to3 = 1'b1;
        end else begin
            ap_idle_pp0_1to3 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage13_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (ap_idle_pp0_0to2 == 1'b1))) begin
            ap_reset_idle_pp0 = 1'b1;
        end else begin
            ap_reset_idle_pp0 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            corners_address0 = zext_ln58_2_fu_1158_p1;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            corners_address0 = zext_ln58_1_fu_1148_p1;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            corners_address0 = zext_ln57_2_fu_1128_p1;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            corners_address0 = zext_ln57_fu_1108_p1;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            corners_address0 = zext_ln56_1_fu_1088_p1;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            corners_address0 = zext_ln55_2_fu_1068_p1;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            corners_address0 = zext_ln55_fu_1048_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            corners_address0 = zext_ln54_1_fu_1028_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            corners_address0 = zext_ln53_2_fu_1008_p1;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            corners_address0 = zext_ln53_fu_988_p1;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            corners_address0 = zext_ln52_1_fu_968_p1;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            corners_address0 = zext_ln51_2_fu_948_p1;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            corners_address0 = zext_ln51_fu_928_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            corners_address0 = zext_ln50_3_fu_655_p1;
        end else begin
            corners_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            corners_address1 = zext_ln58_fu_1138_p1;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            corners_address1 = zext_ln57_1_fu_1118_p1;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            corners_address1 = zext_ln56_2_fu_1098_p1;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            corners_address1 = zext_ln56_fu_1078_p1;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            corners_address1 = zext_ln55_1_fu_1058_p1;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            corners_address1 = zext_ln54_2_fu_1038_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            corners_address1 = zext_ln54_fu_1018_p1;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            corners_address1 = zext_ln53_1_fu_998_p1;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            corners_address1 = zext_ln52_2_fu_978_p1;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            corners_address1 = zext_ln52_fu_958_p1;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            corners_address1 = zext_ln51_1_fu_938_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            corners_address1 = zext_ln50_2_fu_645_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            corners_address1 = zext_ln50_1_fu_544_p1;
        end else begin
            corners_address1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4_11001) 
    & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            corners_ce0 = 1'b1;
        end else begin
            corners_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage1_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            corners_ce1 = 1'b1;
        end else begin
            corners_ce1 = 1'b0;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            corners_d0 = reg_488;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            corners_d0 = reg_494;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            corners_d0 = reg_460;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            corners_d0 = reg_468;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            corners_d0 = add161_2_reg_1418;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            corners_d0 = add6_reg_1413;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            corners_d0 = sub138_1_reg_1408;
        end else if (((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13))) begin
            corners_d0 = reg_500;
        end else if (((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
            corners_d0 = reg_507;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            corners_d0 = reg_524;
        end else if (((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
            corners_d0 = reg_513;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            corners_d0 = tmp_316_fu_764_p6;
        end else begin
            corners_d0 = 'bx;
        end
    end

    always @(*) begin
        if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            corners_d1 = reg_481;
        end else if (((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7))) begin
            corners_d1 = reg_468;
        end else if (((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6))) begin
            corners_d1 = reg_475;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            corners_d1 = reg_460;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            corners_d1 = reg_513;
        end else if ((((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            corners_d1 = reg_529;
        end else if (((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
            corners_d1 = reg_500;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            corners_d1 = reg_519;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            corners_d1 = tmp_315_fu_734_p6;
        end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            corners_d1 = tmp_314_fu_625_p6;
        end else begin
            corners_d1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage9_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4_11001) 
    & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            corners_we0 = 1'b1;
        end else begin
            corners_we0 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage13_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage6_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage1_11001) 
    & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage8_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage7_11001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)))) begin
            corners_we1 = 1'b1;
        end else begin
            corners_we1 = 1'b0;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)))) begin
            grp_fu_419_opcode = 2'd1;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_419_opcode = 2'd0;
        end else begin
            grp_fu_419_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_419_p0 = sub7_reg_1393;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            grp_fu_419_p0 = add5_reg_1378;
        end else if ((((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_419_p0 = sub3_reg_1358;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_419_p0 = reg_500;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_419_p0 = reg_475;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_419_p0 = reg_481;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_419_p0 = reg_460;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_419_p0 = tmp_316_reg_1243_pp0_iter1_reg;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_419_p0 = tmp_314_reg_1216_pp0_iter1_reg;
        end else begin
            grp_fu_419_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_419_p1 = zL_reg_1343_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_419_p1 = zL_reg_1343;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_419_p1 = yL_2_reg_1337;
        end else if ((((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_419_p1 = yL_reg_1326;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_419_p1 = reg_453;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_419_p1 = reg_446;
        end else begin
            grp_fu_419_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
            grp_fu_423_opcode = 2'd1;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_423_opcode = 2'd0;
        end else begin
            grp_fu_423_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_423_p0 = sub204_1_reg_1398;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            grp_fu_423_p0 = add158_1_reg_1383;
        end else if ((((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_423_p0 = sub112_1_reg_1368;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_423_p0 = reg_507;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_423_p0 = reg_488;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)))) begin
            grp_fu_423_p0 = reg_468;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_423_p0 = tmp_315_reg_1238_pp0_iter1_reg;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_423_p0 = tmp_315_reg_1238;
        end else begin
            grp_fu_423_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_423_p1 = zL_1_reg_1348_pp0_iter2_reg;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_423_p1 = zL_1_reg_1348;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_423_p1 = yL_1_reg_1332;
        end else if ((((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_423_p1 = xL_1_reg_1321;
        end else begin
            grp_fu_423_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage0_00001) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage12_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage6_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage4_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage11_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage9_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage2_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage1_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
            grp_fu_427_opcode = 2'd1;
        end else if ((((1'b0 == ap_block_pp0_stage13_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage7_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage5_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage3_00001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage10_00001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_427_opcode = 2'd0;
        end else begin
            grp_fu_427_opcode = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_427_p0 = sub204_2_reg_1403;
        end else if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)))) begin
            grp_fu_427_p0 = add158_2_reg_1388;
        end else if ((((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)))) begin
            grp_fu_427_p0 = sub112_2_reg_1373;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_427_p0 = add67_2_reg_1363;
        end else if ((((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_427_p0 = reg_494;
        end else if (((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
            grp_fu_427_p0 = reg_481;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_427_p0 = reg_460;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_427_p0 = tmp_316_reg_1243_pp0_iter1_reg;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_427_p0 = tmp_314_reg_1216_pp0_iter1_reg;
        end else begin
            grp_fu_427_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage7) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage7)) | ((1'b0 == ap_block_pp0_stage6) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage6)) | ((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5)) | ((1'b0 == ap_block_pp0_stage13) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage13)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
            grp_fu_427_p1 = zL_2_reg_1353_pp0_iter2_reg;
        end else if ((((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4)) | ((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            grp_fu_427_p1 = zL_2_reg_1353;
        end else if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_427_p1 = yL_2_reg_1337;
        end else if (((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
            grp_fu_427_p1 = yL_reg_1326;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_427_p1 = reg_453;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_427_p1 = reg_446;
        end else begin
            grp_fu_427_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage12) & (1'b1 == ap_CS_fsm_pp0_stage12))) begin
                grp_fu_431_p0 = mul1_reg_1316;
            end else if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                grp_fu_431_p0 = mul8_reg_1306;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                grp_fu_431_p0 = mul5_reg_1296;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                grp_fu_431_p0 = reg_453;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                grp_fu_431_p0 = reg_446;
            end else if (((1'b0 == ap_block_pp0_stage5) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
                grp_fu_431_p0 = tmp_313_reg_1281;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                grp_fu_431_p0 = tmp_311_reg_1265;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                grp_fu_431_p0 = tmp_309_reg_1255;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                grp_fu_431_p0 = tmp_307_reg_1228;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                grp_fu_431_p0 = tmp_reg_1206;
            end else begin
                grp_fu_431_p0 = 'bx;
            end
        end else begin
            grp_fu_431_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage12) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage12)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_431_p1 = 64'd4602678819172646912;
        end else if (((1'b0 == ap_block_pp0_stage5) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage5))) begin
            grp_fu_431_p1 = dim_0_2_val_read_reg_1275;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_431_p1 = ap_port_reg_dim_0_2_val;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_431_p1 = dim_0_1_val_read_reg_1249;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_431_p1 = dim_0_0_val_read_reg_1222;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_431_p1 = ap_port_reg_dim_0_0_val;
        end else begin
            grp_fu_431_p1 = 'bx;
        end
    end

    always @(*) begin
        if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
            if (((1'b0 == ap_block_pp0_stage11) & (1'b1 == ap_CS_fsm_pp0_stage11))) begin
                grp_fu_436_p0 = mul9_reg_1311;
            end else if (((1'b0 == ap_block_pp0_stage10) & (1'b1 == ap_CS_fsm_pp0_stage10))) begin
                grp_fu_436_p0 = mul7_reg_1301;
            end else if (((1'b0 == ap_block_pp0_stage9) & (1'b1 == ap_CS_fsm_pp0_stage9))) begin
                grp_fu_436_p0 = mul4_reg_1291;
            end else if (((1'b0 == ap_block_pp0_stage8) & (1'b1 == ap_CS_fsm_pp0_stage8))) begin
                grp_fu_436_p0 = mul6_reg_1286;
            end else if (((1'b0 == ap_block_pp0_stage4) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
                grp_fu_436_p0 = tmp_312_reg_1270;
            end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
                grp_fu_436_p0 = tmp_310_reg_1260;
            end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                grp_fu_436_p0 = tmp_308_reg_1233;
            end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
                grp_fu_436_p0 = tmp_s_reg_1211;
            end else begin
                grp_fu_436_p0 = 'bx;
            end
        end else begin
            grp_fu_436_p0 = 'bx;
        end
    end

    always @(*) begin
        if ((((1'b0 == ap_block_pp0_stage9) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage9)) | ((1'b0 == ap_block_pp0_stage8) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage8)) | ((1'b0 == ap_block_pp0_stage11) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage11)) | ((1'b0 == ap_block_pp0_stage10) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage10)))) begin
            grp_fu_436_p1 = 64'd4602678819172646912;
        end else if (((1'b0 == ap_block_pp0_stage4) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage4))) begin
            grp_fu_436_p1 = ap_port_reg_dim_0_2_val;
        end else if (((1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            grp_fu_436_p1 = dim_0_1_val_read_reg_1249;
        end else if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            grp_fu_436_p1 = ap_port_reg_dim_0_1_val;
        end else if (((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            grp_fu_436_p1 = ap_port_reg_dim_0_0_val;
        end else begin
            grp_fu_436_p1 = 'bx;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_pp0_stage0: begin
                if ((~((ap_start == 1'b0) & (ap_idle_pp0_1to3 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end
            end
            ap_ST_fsm_pp0_stage1: begin
                if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage1;
                end
            end
            ap_ST_fsm_pp0_stage2: begin
                if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage2;
                end
            end
            ap_ST_fsm_pp0_stage3: begin
                if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage3;
                end
            end
            ap_ST_fsm_pp0_stage4: begin
                if ((1'b0 == ap_block_pp0_stage4_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage4;
                end
            end
            ap_ST_fsm_pp0_stage5: begin
                if ((1'b0 == ap_block_pp0_stage5_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage5;
                end
            end
            ap_ST_fsm_pp0_stage6: begin
                if ((1'b0 == ap_block_pp0_stage6_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage6;
                end
            end
            ap_ST_fsm_pp0_stage7: begin
                if ((1'b0 == ap_block_pp0_stage7_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage7;
                end
            end
            ap_ST_fsm_pp0_stage8: begin
                if ((1'b0 == ap_block_pp0_stage8_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage8;
                end
            end
            ap_ST_fsm_pp0_stage9: begin
                if (((1'b0 == ap_block_pp0_stage9_subdone) & (ap_reset_idle_pp0 == 1'b0))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end else if (((1'b0 == ap_block_pp0_stage9_subdone) & (ap_reset_idle_pp0 == 1'b1))) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage9;
                end
            end
            ap_ST_fsm_pp0_stage10: begin
                if ((1'b0 == ap_block_pp0_stage10_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage10;
                end
            end
            ap_ST_fsm_pp0_stage11: begin
                if ((1'b0 == ap_block_pp0_stage11_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage11;
                end
            end
            ap_ST_fsm_pp0_stage12: begin
                if ((1'b0 == ap_block_pp0_stage12_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage12;
                end
            end
            ap_ST_fsm_pp0_stage13: begin
                if ((1'b0 == ap_block_pp0_stage13_subdone)) begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage0;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_pp0_stage13;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign add_ln50_1_fu_650_p2 = (mul_ln50_reg_1176 + 7'd2);

    assign add_ln50_fu_640_p2 = (mul_ln50_reg_1176 + 7'd1);

    assign add_ln51_1_fu_933_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd4);

    assign add_ln51_2_fu_943_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd5);

    assign add_ln51_fu_923_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd3);

    assign add_ln52_1_fu_963_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd7);

    assign add_ln52_2_fu_973_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd8);

    assign add_ln52_fu_953_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd6);

    assign add_ln53_1_fu_993_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd10);

    assign add_ln53_2_fu_1003_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd11);

    assign add_ln53_fu_983_p2 = (mul_ln50_reg_1176_pp0_iter2_reg + 7'd9);

    assign add_ln54_1_fu_1023_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd13);

    assign add_ln54_2_fu_1033_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd14);

    assign add_ln54_fu_1013_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd12);

    assign add_ln55_1_fu_1053_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd16);

    assign add_ln55_2_fu_1063_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd17);

    assign add_ln55_fu_1043_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd15);

    assign add_ln56_1_fu_1083_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd19);

    assign add_ln56_2_fu_1093_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd20);

    assign add_ln56_fu_1073_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd18);

    assign add_ln57_1_fu_1113_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd22);

    assign add_ln57_2_fu_1123_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd23);

    assign add_ln57_fu_1103_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd21);

    assign add_ln58_1_fu_1143_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd25);

    assign add_ln58_2_fu_1153_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd26);

    assign add_ln58_fu_1133_p2 = (mul_ln50_reg_1176_pp0_iter3_reg + 7'd24);

    assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_pp0_stage10 = ap_CS_fsm[32'd10];

    assign ap_CS_fsm_pp0_stage11 = ap_CS_fsm[32'd11];

    assign ap_CS_fsm_pp0_stage12 = ap_CS_fsm[32'd12];

    assign ap_CS_fsm_pp0_stage13 = ap_CS_fsm[32'd13];

    assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd3];

    assign ap_CS_fsm_pp0_stage4 = ap_CS_fsm[32'd4];

    assign ap_CS_fsm_pp0_stage5 = ap_CS_fsm[32'd5];

    assign ap_CS_fsm_pp0_stage6 = ap_CS_fsm[32'd6];

    assign ap_CS_fsm_pp0_stage7 = ap_CS_fsm[32'd7];

    assign ap_CS_fsm_pp0_stage8 = ap_CS_fsm[32'd8];

    assign ap_CS_fsm_pp0_stage9 = ap_CS_fsm[32'd9];

    assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage10_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage11_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage12_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage13_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage4_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage5_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage6_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage7_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage8_subdone = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_00001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_11001 = ~(1'b1 == 1'b1);

    assign ap_block_pp0_stage9_subdone = ~(1'b1 == 1'b1);

    assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

    assign mul_ln50_fu_538_p0 = mul_ln50_fu_538_p00;

    assign mul_ln50_fu_538_p00 = H_offset;

    assign mul_ln50_fu_538_p1 = 7'd27;

    assign zext_ln50_1_fu_544_p1 = mul_ln50_fu_538_p2;

    assign zext_ln50_2_fu_645_p1 = add_ln50_fu_640_p2;

    assign zext_ln50_3_fu_655_p1 = add_ln50_1_fu_650_p2;

    assign zext_ln51_1_fu_938_p1 = add_ln51_1_fu_933_p2;

    assign zext_ln51_2_fu_948_p1 = add_ln51_2_fu_943_p2;

    assign zext_ln51_fu_928_p1 = add_ln51_fu_923_p2;

    assign zext_ln52_1_fu_968_p1 = add_ln52_1_fu_963_p2;

    assign zext_ln52_2_fu_978_p1 = add_ln52_2_fu_973_p2;

    assign zext_ln52_fu_958_p1 = add_ln52_fu_953_p2;

    assign zext_ln53_1_fu_998_p1 = add_ln53_1_fu_993_p2;

    assign zext_ln53_2_fu_1008_p1 = add_ln53_2_fu_1003_p2;

    assign zext_ln53_fu_988_p1 = add_ln53_fu_983_p2;

    assign zext_ln54_1_fu_1028_p1 = add_ln54_1_fu_1023_p2;

    assign zext_ln54_2_fu_1038_p1 = add_ln54_2_fu_1033_p2;

    assign zext_ln54_fu_1018_p1 = add_ln54_fu_1013_p2;

    assign zext_ln55_1_fu_1058_p1 = add_ln55_1_fu_1053_p2;

    assign zext_ln55_2_fu_1068_p1 = add_ln55_2_fu_1063_p2;

    assign zext_ln55_fu_1048_p1 = add_ln55_fu_1043_p2;

    assign zext_ln56_1_fu_1088_p1 = add_ln56_1_fu_1083_p2;

    assign zext_ln56_2_fu_1098_p1 = add_ln56_2_fu_1093_p2;

    assign zext_ln56_fu_1078_p1 = add_ln56_fu_1073_p2;

    assign zext_ln57_1_fu_1118_p1 = add_ln57_1_fu_1113_p2;

    assign zext_ln57_2_fu_1128_p1 = add_ln57_2_fu_1123_p2;

    assign zext_ln57_fu_1108_p1 = add_ln57_fu_1103_p2;

    assign zext_ln58_1_fu_1148_p1 = add_ln58_1_fu_1143_p2;

    assign zext_ln58_2_fu_1158_p1 = add_ln58_2_fu_1153_p2;

    assign zext_ln58_fu_1138_p1 = add_ln58_fu_1133_p2;

endmodule  //main_blockDescToBoundingBox_double_s
