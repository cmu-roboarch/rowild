/*
 * MIT License
 *
 * Copyright (c) 2023 Carnegie Mellon University
 *
 * This file is part of RoWild.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
*/

// ==============================================================
// Generated by Vitis HLS v2023.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// Copyright 2022-2023 Advanced Micro Devices, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module main_forwardKin (
    ap_clk,
    ap_rst,
    ap_start,
    ap_done,
    ap_idle,
    ap_ready,
    this_TLink_0_0_address0,
    this_TLink_0_0_ce0,
    this_TLink_0_0_q0,
    this_TLink_0_1_address0,
    this_TLink_0_1_ce0,
    this_TLink_0_1_q0,
    this_TLink_0_2_address0,
    this_TLink_0_2_ce0,
    this_TLink_0_2_q0,
    this_TLink_0_3_address0,
    this_TLink_0_3_ce0,
    this_TLink_0_3_q0,
    this_TLink_1_0_address0,
    this_TLink_1_0_ce0,
    this_TLink_1_0_q0,
    this_TLink_1_1_address0,
    this_TLink_1_1_ce0,
    this_TLink_1_1_q0,
    this_TLink_1_2_address0,
    this_TLink_1_2_ce0,
    this_TLink_1_2_q0,
    this_TLink_1_3_address0,
    this_TLink_1_3_ce0,
    this_TLink_1_3_q0,
    this_TLink_2_0_address0,
    this_TLink_2_0_ce0,
    this_TLink_2_0_q0,
    this_TLink_2_1_address0,
    this_TLink_2_1_ce0,
    this_TLink_2_1_q0,
    this_TLink_2_2_address0,
    this_TLink_2_2_ce0,
    this_TLink_2_2_q0,
    this_TLink_2_3_address0,
    this_TLink_2_3_ce0,
    this_TLink_2_3_q0,
    this_TLink_3_0_address0,
    this_TLink_3_0_ce0,
    this_TLink_3_0_q0,
    this_TLink_3_1_address0,
    this_TLink_3_1_ce0,
    this_TLink_3_1_q0,
    this_TLink_3_2_address0,
    this_TLink_3_2_ce0,
    this_TLink_3_2_q0,
    this_TLink_3_3_address0,
    this_TLink_3_3_ce0,
    this_TLink_3_3_q0,
    this_TJoint_0_0_address0,
    this_TJoint_0_0_ce0,
    this_TJoint_0_0_we0,
    this_TJoint_0_0_d0,
    this_TJoint_0_0_q0,
    this_TJoint_0_1_address0,
    this_TJoint_0_1_ce0,
    this_TJoint_0_1_we0,
    this_TJoint_0_1_d0,
    this_TJoint_0_1_q0,
    this_TJoint_0_2_address0,
    this_TJoint_0_2_ce0,
    this_TJoint_0_2_we0,
    this_TJoint_0_2_d0,
    this_TJoint_0_2_q0,
    this_TJoint_0_3_address0,
    this_TJoint_0_3_ce0,
    this_TJoint_0_3_we0,
    this_TJoint_0_3_d0,
    this_TJoint_0_3_q0,
    this_TJoint_1_0_address0,
    this_TJoint_1_0_ce0,
    this_TJoint_1_0_we0,
    this_TJoint_1_0_d0,
    this_TJoint_1_0_q0,
    this_TJoint_1_1_address0,
    this_TJoint_1_1_ce0,
    this_TJoint_1_1_we0,
    this_TJoint_1_1_d0,
    this_TJoint_1_1_q0,
    this_TJoint_1_2_address0,
    this_TJoint_1_2_ce0,
    this_TJoint_1_2_we0,
    this_TJoint_1_2_d0,
    this_TJoint_1_2_q0,
    this_TJoint_1_3_address0,
    this_TJoint_1_3_ce0,
    this_TJoint_1_3_we0,
    this_TJoint_1_3_d0,
    this_TJoint_1_3_q0,
    this_TJoint_2_0_address0,
    this_TJoint_2_0_ce0,
    this_TJoint_2_0_we0,
    this_TJoint_2_0_d0,
    this_TJoint_2_0_q0,
    this_TJoint_2_1_address0,
    this_TJoint_2_1_ce0,
    this_TJoint_2_1_we0,
    this_TJoint_2_1_d0,
    this_TJoint_2_1_q0,
    this_TJoint_2_2_address0,
    this_TJoint_2_2_ce0,
    this_TJoint_2_2_we0,
    this_TJoint_2_2_d0,
    this_TJoint_2_2_q0,
    this_TJoint_2_3_address0,
    this_TJoint_2_3_ce0,
    this_TJoint_2_3_we0,
    this_TJoint_2_3_d0,
    this_TJoint_2_3_q0,
    this_TJoint_3_0_address0,
    this_TJoint_3_0_ce0,
    this_TJoint_3_0_we0,
    this_TJoint_3_0_d0,
    this_TJoint_3_0_q0,
    this_TJoint_3_1_address0,
    this_TJoint_3_1_ce0,
    this_TJoint_3_1_we0,
    this_TJoint_3_1_d0,
    this_TJoint_3_1_q0,
    this_TJoint_3_2_address0,
    this_TJoint_3_2_ce0,
    this_TJoint_3_2_we0,
    this_TJoint_3_2_d0,
    this_TJoint_3_2_q0,
    this_TJoint_3_3_address0,
    this_TJoint_3_3_ce0,
    this_TJoint_3_3_we0,
    this_TJoint_3_3_d0,
    this_TJoint_3_3_q0,
    this_TCurr_0_0_address0,
    this_TCurr_0_0_ce0,
    this_TCurr_0_0_we0,
    this_TCurr_0_0_d0,
    this_TCurr_0_0_q0,
    this_TCurr_0_1_address0,
    this_TCurr_0_1_ce0,
    this_TCurr_0_1_we0,
    this_TCurr_0_1_d0,
    this_TCurr_0_1_q0,
    this_TCurr_0_2_address0,
    this_TCurr_0_2_ce0,
    this_TCurr_0_2_we0,
    this_TCurr_0_2_d0,
    this_TCurr_0_2_q0,
    this_TCurr_0_3_address0,
    this_TCurr_0_3_ce0,
    this_TCurr_0_3_we0,
    this_TCurr_0_3_d0,
    this_TCurr_0_3_q0,
    this_TCurr_1_0_address0,
    this_TCurr_1_0_ce0,
    this_TCurr_1_0_we0,
    this_TCurr_1_0_d0,
    this_TCurr_1_0_q0,
    this_TCurr_1_1_address0,
    this_TCurr_1_1_ce0,
    this_TCurr_1_1_we0,
    this_TCurr_1_1_d0,
    this_TCurr_1_1_q0,
    this_TCurr_1_2_address0,
    this_TCurr_1_2_ce0,
    this_TCurr_1_2_we0,
    this_TCurr_1_2_d0,
    this_TCurr_1_2_q0,
    this_TCurr_1_3_address0,
    this_TCurr_1_3_ce0,
    this_TCurr_1_3_we0,
    this_TCurr_1_3_d0,
    this_TCurr_1_3_q0,
    this_TCurr_2_0_address0,
    this_TCurr_2_0_ce0,
    this_TCurr_2_0_we0,
    this_TCurr_2_0_d0,
    this_TCurr_2_0_q0,
    this_TCurr_2_1_address0,
    this_TCurr_2_1_ce0,
    this_TCurr_2_1_we0,
    this_TCurr_2_1_d0,
    this_TCurr_2_1_q0,
    this_TCurr_2_2_address0,
    this_TCurr_2_2_ce0,
    this_TCurr_2_2_we0,
    this_TCurr_2_2_d0,
    this_TCurr_2_2_q0,
    this_TCurr_2_3_address0,
    this_TCurr_2_3_ce0,
    this_TCurr_2_3_we0,
    this_TCurr_2_3_d0,
    this_TCurr_2_3_q0,
    this_TCurr_3_0_address0,
    this_TCurr_3_0_ce0,
    this_TCurr_3_0_we0,
    this_TCurr_3_0_d0,
    this_TCurr_3_0_q0,
    this_TCurr_3_1_address0,
    this_TCurr_3_1_ce0,
    this_TCurr_3_1_we0,
    this_TCurr_3_1_d0,
    this_TCurr_3_1_q0,
    this_TCurr_3_2_address0,
    this_TCurr_3_2_ce0,
    this_TCurr_3_2_we0,
    this_TCurr_3_2_d0,
    this_TCurr_3_2_q0,
    this_TCurr_3_3_address0,
    this_TCurr_3_3_ce0,
    this_TCurr_3_3_we0,
    this_TCurr_3_3_d0,
    this_TCurr_3_3_q0,
    this_q_address0,
    this_q_ce0,
    this_q_we0,
    this_q_d0,
    this_q_q0,
    ang_address0,
    ang_ce0,
    ang_q0
);

    parameter ap_ST_fsm_state1 = 4'd1;
    parameter ap_ST_fsm_state2 = 4'd2;
    parameter ap_ST_fsm_state3 = 4'd4;
    parameter ap_ST_fsm_state4 = 4'd8;

    input ap_clk;
    input ap_rst;
    input ap_start;
    output ap_done;
    output ap_idle;
    output ap_ready;
    output [2:0] this_TLink_0_0_address0;
    output this_TLink_0_0_ce0;
    input [63:0] this_TLink_0_0_q0;
    output [2:0] this_TLink_0_1_address0;
    output this_TLink_0_1_ce0;
    input [63:0] this_TLink_0_1_q0;
    output [2:0] this_TLink_0_2_address0;
    output this_TLink_0_2_ce0;
    input [63:0] this_TLink_0_2_q0;
    output [2:0] this_TLink_0_3_address0;
    output this_TLink_0_3_ce0;
    input [63:0] this_TLink_0_3_q0;
    output [2:0] this_TLink_1_0_address0;
    output this_TLink_1_0_ce0;
    input [63:0] this_TLink_1_0_q0;
    output [2:0] this_TLink_1_1_address0;
    output this_TLink_1_1_ce0;
    input [63:0] this_TLink_1_1_q0;
    output [2:0] this_TLink_1_2_address0;
    output this_TLink_1_2_ce0;
    input [63:0] this_TLink_1_2_q0;
    output [2:0] this_TLink_1_3_address0;
    output this_TLink_1_3_ce0;
    input [63:0] this_TLink_1_3_q0;
    output [2:0] this_TLink_2_0_address0;
    output this_TLink_2_0_ce0;
    input [63:0] this_TLink_2_0_q0;
    output [2:0] this_TLink_2_1_address0;
    output this_TLink_2_1_ce0;
    input [63:0] this_TLink_2_1_q0;
    output [2:0] this_TLink_2_2_address0;
    output this_TLink_2_2_ce0;
    input [63:0] this_TLink_2_2_q0;
    output [2:0] this_TLink_2_3_address0;
    output this_TLink_2_3_ce0;
    input [63:0] this_TLink_2_3_q0;
    output [2:0] this_TLink_3_0_address0;
    output this_TLink_3_0_ce0;
    input [63:0] this_TLink_3_0_q0;
    output [2:0] this_TLink_3_1_address0;
    output this_TLink_3_1_ce0;
    input [63:0] this_TLink_3_1_q0;
    output [2:0] this_TLink_3_2_address0;
    output this_TLink_3_2_ce0;
    input [63:0] this_TLink_3_2_q0;
    output [2:0] this_TLink_3_3_address0;
    output this_TLink_3_3_ce0;
    input [63:0] this_TLink_3_3_q0;
    output [2:0] this_TJoint_0_0_address0;
    output this_TJoint_0_0_ce0;
    output this_TJoint_0_0_we0;
    output [63:0] this_TJoint_0_0_d0;
    input [63:0] this_TJoint_0_0_q0;
    output [2:0] this_TJoint_0_1_address0;
    output this_TJoint_0_1_ce0;
    output this_TJoint_0_1_we0;
    output [63:0] this_TJoint_0_1_d0;
    input [63:0] this_TJoint_0_1_q0;
    output [2:0] this_TJoint_0_2_address0;
    output this_TJoint_0_2_ce0;
    output this_TJoint_0_2_we0;
    output [63:0] this_TJoint_0_2_d0;
    input [63:0] this_TJoint_0_2_q0;
    output [2:0] this_TJoint_0_3_address0;
    output this_TJoint_0_3_ce0;
    output this_TJoint_0_3_we0;
    output [63:0] this_TJoint_0_3_d0;
    input [63:0] this_TJoint_0_3_q0;
    output [2:0] this_TJoint_1_0_address0;
    output this_TJoint_1_0_ce0;
    output this_TJoint_1_0_we0;
    output [63:0] this_TJoint_1_0_d0;
    input [63:0] this_TJoint_1_0_q0;
    output [2:0] this_TJoint_1_1_address0;
    output this_TJoint_1_1_ce0;
    output this_TJoint_1_1_we0;
    output [63:0] this_TJoint_1_1_d0;
    input [63:0] this_TJoint_1_1_q0;
    output [2:0] this_TJoint_1_2_address0;
    output this_TJoint_1_2_ce0;
    output this_TJoint_1_2_we0;
    output [63:0] this_TJoint_1_2_d0;
    input [63:0] this_TJoint_1_2_q0;
    output [2:0] this_TJoint_1_3_address0;
    output this_TJoint_1_3_ce0;
    output this_TJoint_1_3_we0;
    output [63:0] this_TJoint_1_3_d0;
    input [63:0] this_TJoint_1_3_q0;
    output [2:0] this_TJoint_2_0_address0;
    output this_TJoint_2_0_ce0;
    output this_TJoint_2_0_we0;
    output [63:0] this_TJoint_2_0_d0;
    input [63:0] this_TJoint_2_0_q0;
    output [2:0] this_TJoint_2_1_address0;
    output this_TJoint_2_1_ce0;
    output this_TJoint_2_1_we0;
    output [63:0] this_TJoint_2_1_d0;
    input [63:0] this_TJoint_2_1_q0;
    output [2:0] this_TJoint_2_2_address0;
    output this_TJoint_2_2_ce0;
    output this_TJoint_2_2_we0;
    output [63:0] this_TJoint_2_2_d0;
    input [63:0] this_TJoint_2_2_q0;
    output [2:0] this_TJoint_2_3_address0;
    output this_TJoint_2_3_ce0;
    output this_TJoint_2_3_we0;
    output [63:0] this_TJoint_2_3_d0;
    input [63:0] this_TJoint_2_3_q0;
    output [2:0] this_TJoint_3_0_address0;
    output this_TJoint_3_0_ce0;
    output this_TJoint_3_0_we0;
    output [63:0] this_TJoint_3_0_d0;
    input [63:0] this_TJoint_3_0_q0;
    output [2:0] this_TJoint_3_1_address0;
    output this_TJoint_3_1_ce0;
    output this_TJoint_3_1_we0;
    output [63:0] this_TJoint_3_1_d0;
    input [63:0] this_TJoint_3_1_q0;
    output [2:0] this_TJoint_3_2_address0;
    output this_TJoint_3_2_ce0;
    output this_TJoint_3_2_we0;
    output [63:0] this_TJoint_3_2_d0;
    input [63:0] this_TJoint_3_2_q0;
    output [2:0] this_TJoint_3_3_address0;
    output this_TJoint_3_3_ce0;
    output this_TJoint_3_3_we0;
    output [63:0] this_TJoint_3_3_d0;
    input [63:0] this_TJoint_3_3_q0;
    output [2:0] this_TCurr_0_0_address0;
    output this_TCurr_0_0_ce0;
    output this_TCurr_0_0_we0;
    output [63:0] this_TCurr_0_0_d0;
    input [63:0] this_TCurr_0_0_q0;
    output [2:0] this_TCurr_0_1_address0;
    output this_TCurr_0_1_ce0;
    output this_TCurr_0_1_we0;
    output [63:0] this_TCurr_0_1_d0;
    input [63:0] this_TCurr_0_1_q0;
    output [2:0] this_TCurr_0_2_address0;
    output this_TCurr_0_2_ce0;
    output this_TCurr_0_2_we0;
    output [63:0] this_TCurr_0_2_d0;
    input [63:0] this_TCurr_0_2_q0;
    output [2:0] this_TCurr_0_3_address0;
    output this_TCurr_0_3_ce0;
    output this_TCurr_0_3_we0;
    output [63:0] this_TCurr_0_3_d0;
    input [63:0] this_TCurr_0_3_q0;
    output [2:0] this_TCurr_1_0_address0;
    output this_TCurr_1_0_ce0;
    output this_TCurr_1_0_we0;
    output [63:0] this_TCurr_1_0_d0;
    input [63:0] this_TCurr_1_0_q0;
    output [2:0] this_TCurr_1_1_address0;
    output this_TCurr_1_1_ce0;
    output this_TCurr_1_1_we0;
    output [63:0] this_TCurr_1_1_d0;
    input [63:0] this_TCurr_1_1_q0;
    output [2:0] this_TCurr_1_2_address0;
    output this_TCurr_1_2_ce0;
    output this_TCurr_1_2_we0;
    output [63:0] this_TCurr_1_2_d0;
    input [63:0] this_TCurr_1_2_q0;
    output [2:0] this_TCurr_1_3_address0;
    output this_TCurr_1_3_ce0;
    output this_TCurr_1_3_we0;
    output [63:0] this_TCurr_1_3_d0;
    input [63:0] this_TCurr_1_3_q0;
    output [2:0] this_TCurr_2_0_address0;
    output this_TCurr_2_0_ce0;
    output this_TCurr_2_0_we0;
    output [63:0] this_TCurr_2_0_d0;
    input [63:0] this_TCurr_2_0_q0;
    output [2:0] this_TCurr_2_1_address0;
    output this_TCurr_2_1_ce0;
    output this_TCurr_2_1_we0;
    output [63:0] this_TCurr_2_1_d0;
    input [63:0] this_TCurr_2_1_q0;
    output [2:0] this_TCurr_2_2_address0;
    output this_TCurr_2_2_ce0;
    output this_TCurr_2_2_we0;
    output [63:0] this_TCurr_2_2_d0;
    input [63:0] this_TCurr_2_2_q0;
    output [2:0] this_TCurr_2_3_address0;
    output this_TCurr_2_3_ce0;
    output this_TCurr_2_3_we0;
    output [63:0] this_TCurr_2_3_d0;
    input [63:0] this_TCurr_2_3_q0;
    output [2:0] this_TCurr_3_0_address0;
    output this_TCurr_3_0_ce0;
    output this_TCurr_3_0_we0;
    output [63:0] this_TCurr_3_0_d0;
    input [63:0] this_TCurr_3_0_q0;
    output [2:0] this_TCurr_3_1_address0;
    output this_TCurr_3_1_ce0;
    output this_TCurr_3_1_we0;
    output [63:0] this_TCurr_3_1_d0;
    input [63:0] this_TCurr_3_1_q0;
    output [2:0] this_TCurr_3_2_address0;
    output this_TCurr_3_2_ce0;
    output this_TCurr_3_2_we0;
    output [63:0] this_TCurr_3_2_d0;
    input [63:0] this_TCurr_3_2_q0;
    output [2:0] this_TCurr_3_3_address0;
    output this_TCurr_3_3_ce0;
    output this_TCurr_3_3_we0;
    output [63:0] this_TCurr_3_3_d0;
    input [63:0] this_TCurr_3_3_q0;
    output [2:0] this_q_address0;
    output this_q_ce0;
    output this_q_we0;
    output [63:0] this_q_d0;
    input [63:0] this_q_q0;
    output [2:0] ang_address0;
    output ang_ce0;
    input [63:0] ang_q0;

    reg ap_done;
    reg ap_idle;
    reg ap_ready;
    reg[2:0] this_TLink_0_0_address0;
    reg this_TLink_0_0_ce0;
    reg[2:0] this_TLink_0_1_address0;
    reg this_TLink_0_1_ce0;
    reg[2:0] this_TLink_0_2_address0;
    reg this_TLink_0_2_ce0;
    reg[2:0] this_TLink_0_3_address0;
    reg this_TLink_0_3_ce0;
    reg[2:0] this_TLink_1_0_address0;
    reg this_TLink_1_0_ce0;
    reg[2:0] this_TLink_1_1_address0;
    reg this_TLink_1_1_ce0;
    reg[2:0] this_TLink_1_2_address0;
    reg this_TLink_1_2_ce0;
    reg[2:0] this_TLink_1_3_address0;
    reg this_TLink_1_3_ce0;
    reg[2:0] this_TLink_2_0_address0;
    reg this_TLink_2_0_ce0;
    reg[2:0] this_TLink_2_1_address0;
    reg this_TLink_2_1_ce0;
    reg[2:0] this_TLink_2_2_address0;
    reg this_TLink_2_2_ce0;
    reg[2:0] this_TLink_2_3_address0;
    reg this_TLink_2_3_ce0;
    reg[2:0] this_TLink_3_0_address0;
    reg this_TLink_3_0_ce0;
    reg[2:0] this_TLink_3_1_address0;
    reg this_TLink_3_1_ce0;
    reg[2:0] this_TLink_3_2_address0;
    reg this_TLink_3_2_ce0;
    reg[2:0] this_TLink_3_3_address0;
    reg this_TLink_3_3_ce0;
    reg[2:0] this_q_address0;
    reg this_q_ce0;
    reg this_q_we0;

    (* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
    wire    ap_CS_fsm_state1;
    reg   [63:0] this_TLink_0_0_load_reg_572;
    wire    ap_CS_fsm_state2;
    reg   [63:0] this_TLink_0_1_load_reg_577;
    reg   [63:0] this_TLink_0_2_load_reg_582;
    reg   [63:0] this_TLink_0_3_load_reg_587;
    reg   [63:0] this_TLink_1_0_load_reg_592;
    reg   [63:0] this_TLink_1_1_load_reg_597;
    reg   [63:0] this_TLink_1_2_load_reg_602;
    reg   [63:0] this_TLink_1_3_load_reg_607;
    reg   [63:0] this_TLink_2_0_load_reg_612;
    reg   [63:0] this_TLink_2_1_load_reg_617;
    reg   [63:0] this_TLink_2_2_load_reg_622;
    reg   [63:0] this_TLink_2_3_load_reg_627;
    reg   [63:0] this_TLink_3_0_load_reg_632;
    reg   [63:0] this_TLink_3_1_load_reg_637;
    reg   [63:0] this_TLink_3_2_load_reg_642;
    reg   [63:0] this_TLink_3_3_load_reg_647;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_done;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_idle;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_ready;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_d0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_idle;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_ready;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_ce0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_we0;
    wire   [63:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_d0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_ce0;
    wire   [2:0] grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_address0;
    wire    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_ce0;
    reg    grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg;
    reg    grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg;
    wire    ap_CS_fsm_state3;
    wire    ap_CS_fsm_state4;
    reg   [3:0] ap_NS_fsm;
    reg    ap_ST_fsm_state1_blk;
    reg    ap_ST_fsm_state2_blk;
    wire    ap_ST_fsm_state3_blk;
    reg    ap_ST_fsm_state4_blk;
    wire    ap_ce_reg;

    // power-on initialization
    initial begin
        #0 ap_CS_fsm = 4'd1;
        #0 grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg = 1'b0;
        #0 grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg = 1'b0;
    end

    main_forwardKin_Pipeline_VITIS_LOOP_202_1 grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start),
        .ap_done(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_done),
        .ap_idle(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_idle),
        .ap_ready(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_ready),
        .ang_address0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_address0),
        .ang_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_ce0),
        .ang_q0(ang_q0),
        .this_q_address0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_address0),
        .this_q_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_ce0),
        .this_q_we0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_we0),
        .this_q_d0(grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_d0)
    );

    main_forwardKin_Pipeline_VITIS_LOOP_218_3 grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356 (
        .ap_clk(ap_clk),
        .ap_rst(ap_rst),
        .ap_start(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start),
        .ap_done(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done),
        .ap_idle(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_idle),
        .ap_ready(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_ready),
        .this_TLink_0_0_load(this_TLink_0_0_load_reg_572),
        .this_TLink_0_1_load(this_TLink_0_1_load_reg_577),
        .this_TLink_0_2_load(this_TLink_0_2_load_reg_582),
        .this_TLink_0_3_load(this_TLink_0_3_load_reg_587),
        .this_TLink_1_0_load(this_TLink_1_0_load_reg_592),
        .this_TLink_1_1_load(this_TLink_1_1_load_reg_597),
        .this_TLink_1_2_load(this_TLink_1_2_load_reg_602),
        .this_TLink_1_3_load(this_TLink_1_3_load_reg_607),
        .this_TLink_2_0_load(this_TLink_2_0_load_reg_612),
        .this_TLink_2_1_load(this_TLink_2_1_load_reg_617),
        .this_TLink_2_2_load(this_TLink_2_2_load_reg_622),
        .this_TLink_2_3_load(this_TLink_2_3_load_reg_627),
        .this_TLink_3_0_load(this_TLink_3_0_load_reg_632),
        .this_TLink_3_1_load(this_TLink_3_1_load_reg_637),
        .this_TLink_3_2_load(this_TLink_3_2_load_reg_642),
        .this_TLink_3_3_load(this_TLink_3_3_load_reg_647),
        .this_TJoint_0_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_address0),
        .this_TJoint_0_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_ce0),
        .this_TJoint_0_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_we0),
        .this_TJoint_0_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_d0),
        .this_TJoint_0_0_q0(this_TJoint_0_0_q0),
        .this_TJoint_1_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_address0),
        .this_TJoint_1_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_ce0),
        .this_TJoint_1_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_we0),
        .this_TJoint_1_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_d0),
        .this_TJoint_1_0_q0(this_TJoint_1_0_q0),
        .this_TJoint_2_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_address0),
        .this_TJoint_2_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_ce0),
        .this_TJoint_2_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_we0),
        .this_TJoint_2_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_d0),
        .this_TJoint_2_0_q0(this_TJoint_2_0_q0),
        .this_TJoint_3_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_address0),
        .this_TJoint_3_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_ce0),
        .this_TJoint_3_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_we0),
        .this_TJoint_3_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_d0),
        .this_TJoint_3_0_q0(this_TJoint_3_0_q0),
        .this_TCurr_0_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_address0),
        .this_TCurr_0_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_ce0),
        .this_TCurr_0_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_we0),
        .this_TCurr_0_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_d0),
        .this_TCurr_0_0_q0(this_TCurr_0_0_q0),
        .this_TJoint_0_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_address0),
        .this_TJoint_0_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_ce0),
        .this_TJoint_0_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_we0),
        .this_TJoint_0_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_d0),
        .this_TJoint_0_1_q0(this_TJoint_0_1_q0),
        .this_TJoint_1_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_address0),
        .this_TJoint_1_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_ce0),
        .this_TJoint_1_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_we0),
        .this_TJoint_1_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_d0),
        .this_TJoint_1_1_q0(this_TJoint_1_1_q0),
        .this_TJoint_2_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_address0),
        .this_TJoint_2_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_ce0),
        .this_TJoint_2_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_we0),
        .this_TJoint_2_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_d0),
        .this_TJoint_2_1_q0(this_TJoint_2_1_q0),
        .this_TJoint_3_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_address0),
        .this_TJoint_3_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_ce0),
        .this_TJoint_3_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_we0),
        .this_TJoint_3_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_d0),
        .this_TJoint_3_1_q0(this_TJoint_3_1_q0),
        .this_TCurr_0_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_address0),
        .this_TCurr_0_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_ce0),
        .this_TCurr_0_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_we0),
        .this_TCurr_0_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_d0),
        .this_TCurr_0_1_q0(this_TCurr_0_1_q0),
        .this_TJoint_0_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_address0),
        .this_TJoint_0_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_ce0),
        .this_TJoint_0_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_we0),
        .this_TJoint_0_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_d0),
        .this_TJoint_0_2_q0(this_TJoint_0_2_q0),
        .this_TJoint_1_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_address0),
        .this_TJoint_1_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_ce0),
        .this_TJoint_1_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_we0),
        .this_TJoint_1_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_d0),
        .this_TJoint_1_2_q0(this_TJoint_1_2_q0),
        .this_TJoint_2_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_address0),
        .this_TJoint_2_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_ce0),
        .this_TJoint_2_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_we0),
        .this_TJoint_2_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_d0),
        .this_TJoint_2_2_q0(this_TJoint_2_2_q0),
        .this_TJoint_3_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_address0),
        .this_TJoint_3_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_ce0),
        .this_TJoint_3_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_we0),
        .this_TJoint_3_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_d0),
        .this_TJoint_3_2_q0(this_TJoint_3_2_q0),
        .this_TCurr_0_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_address0),
        .this_TCurr_0_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_ce0),
        .this_TCurr_0_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_we0),
        .this_TCurr_0_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_d0),
        .this_TCurr_0_2_q0(this_TCurr_0_2_q0),
        .this_TJoint_0_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_address0),
        .this_TJoint_0_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_ce0),
        .this_TJoint_0_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_we0),
        .this_TJoint_0_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_d0),
        .this_TJoint_0_3_q0(this_TJoint_0_3_q0),
        .this_TJoint_1_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_address0),
        .this_TJoint_1_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_ce0),
        .this_TJoint_1_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_we0),
        .this_TJoint_1_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_d0),
        .this_TJoint_1_3_q0(this_TJoint_1_3_q0),
        .this_TJoint_2_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_address0),
        .this_TJoint_2_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_ce0),
        .this_TJoint_2_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_we0),
        .this_TJoint_2_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_d0),
        .this_TJoint_2_3_q0(this_TJoint_2_3_q0),
        .this_TJoint_3_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_address0),
        .this_TJoint_3_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_ce0),
        .this_TJoint_3_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_we0),
        .this_TJoint_3_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_d0),
        .this_TJoint_3_3_q0(this_TJoint_3_3_q0),
        .this_TCurr_0_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_address0),
        .this_TCurr_0_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_ce0),
        .this_TCurr_0_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_we0),
        .this_TCurr_0_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_d0),
        .this_TCurr_0_3_q0(this_TCurr_0_3_q0),
        .this_TCurr_1_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_address0),
        .this_TCurr_1_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_ce0),
        .this_TCurr_1_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_we0),
        .this_TCurr_1_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_d0),
        .this_TCurr_1_0_q0(this_TCurr_1_0_q0),
        .this_TCurr_1_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_address0),
        .this_TCurr_1_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_ce0),
        .this_TCurr_1_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_we0),
        .this_TCurr_1_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_d0),
        .this_TCurr_1_1_q0(this_TCurr_1_1_q0),
        .this_TCurr_1_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_address0),
        .this_TCurr_1_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_ce0),
        .this_TCurr_1_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_we0),
        .this_TCurr_1_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_d0),
        .this_TCurr_1_2_q0(this_TCurr_1_2_q0),
        .this_TCurr_1_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_address0),
        .this_TCurr_1_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_ce0),
        .this_TCurr_1_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_we0),
        .this_TCurr_1_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_d0),
        .this_TCurr_1_3_q0(this_TCurr_1_3_q0),
        .this_TCurr_2_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_address0),
        .this_TCurr_2_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_ce0),
        .this_TCurr_2_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_we0),
        .this_TCurr_2_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_d0),
        .this_TCurr_2_0_q0(this_TCurr_2_0_q0),
        .this_TCurr_2_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_address0),
        .this_TCurr_2_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_ce0),
        .this_TCurr_2_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_we0),
        .this_TCurr_2_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_d0),
        .this_TCurr_2_1_q0(this_TCurr_2_1_q0),
        .this_TCurr_2_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_address0),
        .this_TCurr_2_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_ce0),
        .this_TCurr_2_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_we0),
        .this_TCurr_2_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_d0),
        .this_TCurr_2_2_q0(this_TCurr_2_2_q0),
        .this_TCurr_2_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_address0),
        .this_TCurr_2_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_ce0),
        .this_TCurr_2_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_we0),
        .this_TCurr_2_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_d0),
        .this_TCurr_2_3_q0(this_TCurr_2_3_q0),
        .this_TCurr_3_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_address0),
        .this_TCurr_3_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_ce0),
        .this_TCurr_3_0_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_we0),
        .this_TCurr_3_0_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_d0),
        .this_TCurr_3_0_q0(this_TCurr_3_0_q0),
        .this_TCurr_3_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_address0),
        .this_TCurr_3_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_ce0),
        .this_TCurr_3_1_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_we0),
        .this_TCurr_3_1_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_d0),
        .this_TCurr_3_1_q0(this_TCurr_3_1_q0),
        .this_TCurr_3_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_address0),
        .this_TCurr_3_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_ce0),
        .this_TCurr_3_2_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_we0),
        .this_TCurr_3_2_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_d0),
        .this_TCurr_3_2_q0(this_TCurr_3_2_q0),
        .this_TCurr_3_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_address0),
        .this_TCurr_3_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_ce0),
        .this_TCurr_3_3_we0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_we0),
        .this_TCurr_3_3_d0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_d0),
        .this_TCurr_3_3_q0(this_TCurr_3_3_q0),
        .this_q_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_address0),
        .this_q_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_ce0),
        .this_q_q0(this_q_q0),
        .this_TLink_0_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_address0),
        .this_TLink_0_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_ce0),
        .this_TLink_0_0_q0(this_TLink_0_0_q0),
        .this_TLink_1_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_address0),
        .this_TLink_1_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_ce0),
        .this_TLink_1_0_q0(this_TLink_1_0_q0),
        .this_TLink_2_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_address0),
        .this_TLink_2_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_ce0),
        .this_TLink_2_0_q0(this_TLink_2_0_q0),
        .this_TLink_3_0_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_address0),
        .this_TLink_3_0_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_ce0),
        .this_TLink_3_0_q0(this_TLink_3_0_q0),
        .this_TLink_0_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_address0),
        .this_TLink_0_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_ce0),
        .this_TLink_0_1_q0(this_TLink_0_1_q0),
        .this_TLink_1_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_address0),
        .this_TLink_1_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_ce0),
        .this_TLink_1_1_q0(this_TLink_1_1_q0),
        .this_TLink_2_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_address0),
        .this_TLink_2_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_ce0),
        .this_TLink_2_1_q0(this_TLink_2_1_q0),
        .this_TLink_3_1_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_address0),
        .this_TLink_3_1_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_ce0),
        .this_TLink_3_1_q0(this_TLink_3_1_q0),
        .this_TLink_0_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_address0),
        .this_TLink_0_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_ce0),
        .this_TLink_0_2_q0(this_TLink_0_2_q0),
        .this_TLink_1_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_address0),
        .this_TLink_1_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_ce0),
        .this_TLink_1_2_q0(this_TLink_1_2_q0),
        .this_TLink_2_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_address0),
        .this_TLink_2_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_ce0),
        .this_TLink_2_2_q0(this_TLink_2_2_q0),
        .this_TLink_3_2_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_address0),
        .this_TLink_3_2_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_ce0),
        .this_TLink_3_2_q0(this_TLink_3_2_q0),
        .this_TLink_0_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_address0),
        .this_TLink_0_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_ce0),
        .this_TLink_0_3_q0(this_TLink_0_3_q0),
        .this_TLink_1_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_address0),
        .this_TLink_1_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_ce0),
        .this_TLink_1_3_q0(this_TLink_1_3_q0),
        .this_TLink_2_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_address0),
        .this_TLink_2_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_ce0),
        .this_TLink_2_3_q0(this_TLink_2_3_q0),
        .this_TLink_3_3_address0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_address0),
        .this_TLink_3_3_ce0(grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_ce0),
        .this_TLink_3_3_q0(this_TLink_3_3_q0)
    );

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            ap_CS_fsm <= ap_ST_fsm_state1;
        end else begin
            ap_CS_fsm <= ap_NS_fsm;
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg <= 1'b0;
        end else begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg <= 1'b1;
            end else if ((grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_ready == 1'b1)) begin
                grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if (ap_rst == 1'b1) begin
            grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg <= 1'b0;
        end else begin
            if ((1'b1 == ap_CS_fsm_state3)) begin
                grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg <= 1'b1;
            end else if ((grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_ready == 1'b1)) begin
                grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg <= 1'b0;
            end
        end
    end

    always @(posedge ap_clk) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_TLink_0_0_load_reg_572 <= this_TLink_0_0_q0;
            this_TLink_0_1_load_reg_577 <= this_TLink_0_1_q0;
            this_TLink_0_2_load_reg_582 <= this_TLink_0_2_q0;
            this_TLink_0_3_load_reg_587 <= this_TLink_0_3_q0;
            this_TLink_1_0_load_reg_592 <= this_TLink_1_0_q0;
            this_TLink_1_1_load_reg_597 <= this_TLink_1_1_q0;
            this_TLink_1_2_load_reg_602 <= this_TLink_1_2_q0;
            this_TLink_1_3_load_reg_607 <= this_TLink_1_3_q0;
            this_TLink_2_0_load_reg_612 <= this_TLink_2_0_q0;
            this_TLink_2_1_load_reg_617 <= this_TLink_2_1_q0;
            this_TLink_2_2_load_reg_622 <= this_TLink_2_2_q0;
            this_TLink_2_3_load_reg_627 <= this_TLink_2_3_q0;
            this_TLink_3_0_load_reg_632 <= this_TLink_3_0_q0;
            this_TLink_3_1_load_reg_637 <= this_TLink_3_1_q0;
            this_TLink_3_2_load_reg_642 <= this_TLink_3_2_q0;
            this_TLink_3_3_load_reg_647 <= this_TLink_3_3_q0;
        end
    end

    always @(*) begin
        if ((ap_start == 1'b0)) begin
            ap_ST_fsm_state1_blk = 1'b1;
        end else begin
            ap_ST_fsm_state1_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_done == 1'b0)) begin
            ap_ST_fsm_state2_blk = 1'b1;
        end else begin
            ap_ST_fsm_state2_blk = 1'b0;
        end
    end

    assign ap_ST_fsm_state3_blk = 1'b0;

    always @(*) begin
        if ((grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done == 1'b0)) begin
            ap_ST_fsm_state4_blk = 1'b1;
        end else begin
            ap_ST_fsm_state4_blk = 1'b0;
        end
    end

    always @(*) begin
        if ((((grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state4)) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_done = 1'b1;
        end else begin
            ap_done = 1'b0;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_idle = 1'b1;
        end else begin
            ap_idle = 1'b0;
        end
    end

    always @(*) begin
        if (((grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state4))) begin
            ap_ready = 1'b1;
        end else begin
            ap_ready = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_0_0_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_address0;
        end else begin
            this_TLink_0_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_0_0_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_0_ce0;
        end else begin
            this_TLink_0_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_0_1_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_address0;
        end else begin
            this_TLink_0_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_0_1_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_1_ce0;
        end else begin
            this_TLink_0_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_0_2_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_address0;
        end else begin
            this_TLink_0_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_0_2_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_2_ce0;
        end else begin
            this_TLink_0_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_0_3_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_address0;
        end else begin
            this_TLink_0_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_0_3_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_0_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_0_3_ce0;
        end else begin
            this_TLink_0_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_1_0_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_address0;
        end else begin
            this_TLink_1_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_1_0_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_0_ce0;
        end else begin
            this_TLink_1_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_1_1_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_address0;
        end else begin
            this_TLink_1_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_1_1_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_1_ce0;
        end else begin
            this_TLink_1_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_1_2_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_address0;
        end else begin
            this_TLink_1_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_1_2_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_2_ce0;
        end else begin
            this_TLink_1_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_1_3_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_address0;
        end else begin
            this_TLink_1_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_1_3_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_1_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_1_3_ce0;
        end else begin
            this_TLink_1_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_2_0_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_address0;
        end else begin
            this_TLink_2_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_2_0_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_0_ce0;
        end else begin
            this_TLink_2_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_2_1_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_address0;
        end else begin
            this_TLink_2_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_2_1_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_1_ce0;
        end else begin
            this_TLink_2_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_2_2_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_address0;
        end else begin
            this_TLink_2_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_2_2_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_2_ce0;
        end else begin
            this_TLink_2_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_2_3_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_address0;
        end else begin
            this_TLink_2_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_2_3_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_2_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_2_3_ce0;
        end else begin
            this_TLink_2_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_3_0_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_address0;
        end else begin
            this_TLink_3_0_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_3_0_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_0_ce0;
        end else begin
            this_TLink_3_0_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_3_1_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_address0;
        end else begin
            this_TLink_3_1_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_3_1_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_1_ce0;
        end else begin
            this_TLink_3_1_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_3_2_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_address0;
        end else begin
            this_TLink_3_2_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_3_2_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_2_ce0;
        end else begin
            this_TLink_3_2_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state1)) begin
            this_TLink_3_3_address0 = 64'd0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_address0;
        end else begin
            this_TLink_3_3_address0 = 'bx;
        end
    end

    always @(*) begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            this_TLink_3_3_ce0 = 1'b1;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            this_TLink_3_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TLink_3_3_ce0;
        end else begin
            this_TLink_3_3_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_q_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_address0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_q_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_address0;
        end else begin
            this_q_address0 = 'bx;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state4)) begin
            this_q_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_q_ce0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            this_q_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_ce0;
        end else begin
            this_q_ce0 = 1'b0;
        end
    end

    always @(*) begin
        if ((1'b1 == ap_CS_fsm_state2)) begin
            this_q_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_we0;
        end else begin
            this_q_we0 = 1'b0;
        end
    end

    always @(*) begin
        case (ap_CS_fsm)
            ap_ST_fsm_state1: begin
                if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end
            end
            ap_ST_fsm_state2: begin
                if (((grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state2))) begin
                    ap_NS_fsm = ap_ST_fsm_state3;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state2;
                end
            end
            ap_ST_fsm_state3: begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
            ap_ST_fsm_state4: begin
                if (((grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state4))) begin
                    ap_NS_fsm = ap_ST_fsm_state1;
                end else begin
                    ap_NS_fsm = ap_ST_fsm_state4;
                end
            end
            default: begin
                ap_NS_fsm = 'bx;
            end
        endcase
    end

    assign ang_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_address0;

    assign ang_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ang_ce0;

    assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

    assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

    assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

    assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

    assign grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_ap_start_reg;

    assign grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_ap_start_reg;

    assign this_TCurr_0_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_address0;

    assign this_TCurr_0_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_ce0;

    assign this_TCurr_0_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_d0;

    assign this_TCurr_0_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_0_we0;

    assign this_TCurr_0_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_address0;

    assign this_TCurr_0_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_ce0;

    assign this_TCurr_0_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_d0;

    assign this_TCurr_0_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_1_we0;

    assign this_TCurr_0_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_address0;

    assign this_TCurr_0_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_ce0;

    assign this_TCurr_0_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_d0;

    assign this_TCurr_0_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_2_we0;

    assign this_TCurr_0_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_address0;

    assign this_TCurr_0_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_ce0;

    assign this_TCurr_0_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_d0;

    assign this_TCurr_0_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_0_3_we0;

    assign this_TCurr_1_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_address0;

    assign this_TCurr_1_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_ce0;

    assign this_TCurr_1_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_d0;

    assign this_TCurr_1_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_0_we0;

    assign this_TCurr_1_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_address0;

    assign this_TCurr_1_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_ce0;

    assign this_TCurr_1_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_d0;

    assign this_TCurr_1_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_1_we0;

    assign this_TCurr_1_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_address0;

    assign this_TCurr_1_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_ce0;

    assign this_TCurr_1_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_d0;

    assign this_TCurr_1_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_2_we0;

    assign this_TCurr_1_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_address0;

    assign this_TCurr_1_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_ce0;

    assign this_TCurr_1_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_d0;

    assign this_TCurr_1_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_1_3_we0;

    assign this_TCurr_2_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_address0;

    assign this_TCurr_2_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_ce0;

    assign this_TCurr_2_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_d0;

    assign this_TCurr_2_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_0_we0;

    assign this_TCurr_2_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_address0;

    assign this_TCurr_2_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_ce0;

    assign this_TCurr_2_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_d0;

    assign this_TCurr_2_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_1_we0;

    assign this_TCurr_2_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_address0;

    assign this_TCurr_2_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_ce0;

    assign this_TCurr_2_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_d0;

    assign this_TCurr_2_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_2_we0;

    assign this_TCurr_2_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_address0;

    assign this_TCurr_2_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_ce0;

    assign this_TCurr_2_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_d0;

    assign this_TCurr_2_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_2_3_we0;

    assign this_TCurr_3_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_address0;

    assign this_TCurr_3_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_ce0;

    assign this_TCurr_3_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_d0;

    assign this_TCurr_3_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_0_we0;

    assign this_TCurr_3_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_address0;

    assign this_TCurr_3_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_ce0;

    assign this_TCurr_3_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_d0;

    assign this_TCurr_3_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_1_we0;

    assign this_TCurr_3_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_address0;

    assign this_TCurr_3_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_ce0;

    assign this_TCurr_3_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_d0;

    assign this_TCurr_3_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_2_we0;

    assign this_TCurr_3_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_address0;

    assign this_TCurr_3_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_ce0;

    assign this_TCurr_3_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_d0;

    assign this_TCurr_3_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TCurr_3_3_we0;

    assign this_TJoint_0_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_address0;

    assign this_TJoint_0_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_ce0;

    assign this_TJoint_0_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_d0;

    assign this_TJoint_0_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_0_we0;

    assign this_TJoint_0_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_address0;

    assign this_TJoint_0_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_ce0;

    assign this_TJoint_0_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_d0;

    assign this_TJoint_0_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_1_we0;

    assign this_TJoint_0_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_address0;

    assign this_TJoint_0_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_ce0;

    assign this_TJoint_0_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_d0;

    assign this_TJoint_0_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_2_we0;

    assign this_TJoint_0_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_address0;

    assign this_TJoint_0_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_ce0;

    assign this_TJoint_0_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_d0;

    assign this_TJoint_0_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_0_3_we0;

    assign this_TJoint_1_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_address0;

    assign this_TJoint_1_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_ce0;

    assign this_TJoint_1_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_d0;

    assign this_TJoint_1_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_0_we0;

    assign this_TJoint_1_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_address0;

    assign this_TJoint_1_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_ce0;

    assign this_TJoint_1_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_d0;

    assign this_TJoint_1_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_1_we0;

    assign this_TJoint_1_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_address0;

    assign this_TJoint_1_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_ce0;

    assign this_TJoint_1_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_d0;

    assign this_TJoint_1_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_2_we0;

    assign this_TJoint_1_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_address0;

    assign this_TJoint_1_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_ce0;

    assign this_TJoint_1_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_d0;

    assign this_TJoint_1_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_1_3_we0;

    assign this_TJoint_2_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_address0;

    assign this_TJoint_2_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_ce0;

    assign this_TJoint_2_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_d0;

    assign this_TJoint_2_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_0_we0;

    assign this_TJoint_2_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_address0;

    assign this_TJoint_2_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_ce0;

    assign this_TJoint_2_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_d0;

    assign this_TJoint_2_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_1_we0;

    assign this_TJoint_2_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_address0;

    assign this_TJoint_2_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_ce0;

    assign this_TJoint_2_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_d0;

    assign this_TJoint_2_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_2_we0;

    assign this_TJoint_2_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_address0;

    assign this_TJoint_2_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_ce0;

    assign this_TJoint_2_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_d0;

    assign this_TJoint_2_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_2_3_we0;

    assign this_TJoint_3_0_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_address0;

    assign this_TJoint_3_0_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_ce0;

    assign this_TJoint_3_0_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_d0;

    assign this_TJoint_3_0_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_0_we0;

    assign this_TJoint_3_1_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_address0;

    assign this_TJoint_3_1_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_ce0;

    assign this_TJoint_3_1_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_d0;

    assign this_TJoint_3_1_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_1_we0;

    assign this_TJoint_3_2_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_address0;

    assign this_TJoint_3_2_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_ce0;

    assign this_TJoint_3_2_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_d0;

    assign this_TJoint_3_2_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_2_we0;

    assign this_TJoint_3_3_address0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_address0;

    assign this_TJoint_3_3_ce0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_ce0;

    assign this_TJoint_3_3_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_d0;

    assign this_TJoint_3_3_we0 = grp_forwardKin_Pipeline_VITIS_LOOP_218_3_fu_356_this_TJoint_3_3_we0;

    assign this_q_d0 = grp_forwardKin_Pipeline_VITIS_LOOP_202_1_fu_348_this_q_d0;

endmodule  //main_forwardKin
